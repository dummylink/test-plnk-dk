--megafunction wizard: %Altera SOPC Builder%
--GENERATION: STANDARD
--VERSION: WM1.0


--Legal Notice: (C)2010 Altera Corporation. All rights reserved.  Your
--use of Altera Corporation's design tools, logic functions and other
--software and tools, and its AMPP partner logic functions, and any
--output files any of the foregoing (including device programming or
--simulation files), and any associated documentation or information are
--expressly subject to the terms and conditions of the Altera Program
--License Subscription Agreement or other applicable license agreement,
--including, without limitation, that your use is for the sole purpose
--of programming logic devices manufactured by Altera and sold by Altera
--or its authorized distributors.  Please refer to the applicable
--agreement for further details.


-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity OpenMAC_0_CMP_arbitrator is 
        port (
              -- inputs:
                 signal OpenMAC_0_CMP_irq : IN STD_LOGIC;
                 signal OpenMAC_0_CMP_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal clk : IN STD_LOGIC;
                 signal niosII_openMac_clock_1_out_address_to_slave : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal niosII_openMac_clock_1_out_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal niosII_openMac_clock_1_out_read : IN STD_LOGIC;
                 signal niosII_openMac_clock_1_out_write : IN STD_LOGIC;
                 signal niosII_openMac_clock_1_out_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal OpenMAC_0_CMP_address : OUT STD_LOGIC;
                 signal OpenMAC_0_CMP_byteenable_n : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal OpenMAC_0_CMP_chipselect : OUT STD_LOGIC;
                 signal OpenMAC_0_CMP_irq_from_sa : OUT STD_LOGIC;
                 signal OpenMAC_0_CMP_read_n : OUT STD_LOGIC;
                 signal OpenMAC_0_CMP_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal OpenMAC_0_CMP_reset_n : OUT STD_LOGIC;
                 signal OpenMAC_0_CMP_write_n : OUT STD_LOGIC;
                 signal OpenMAC_0_CMP_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal d1_OpenMAC_0_CMP_end_xfer : OUT STD_LOGIC;
                 signal niosII_openMac_clock_1_out_granted_OpenMAC_0_CMP : OUT STD_LOGIC;
                 signal niosII_openMac_clock_1_out_qualified_request_OpenMAC_0_CMP : OUT STD_LOGIC;
                 signal niosII_openMac_clock_1_out_read_data_valid_OpenMAC_0_CMP : OUT STD_LOGIC;
                 signal niosII_openMac_clock_1_out_requests_OpenMAC_0_CMP : OUT STD_LOGIC
              );
end entity OpenMAC_0_CMP_arbitrator;


architecture europa of OpenMAC_0_CMP_arbitrator is
                signal OpenMAC_0_CMP_allgrants :  STD_LOGIC;
                signal OpenMAC_0_CMP_allow_new_arb_cycle :  STD_LOGIC;
                signal OpenMAC_0_CMP_any_bursting_master_saved_grant :  STD_LOGIC;
                signal OpenMAC_0_CMP_any_continuerequest :  STD_LOGIC;
                signal OpenMAC_0_CMP_arb_counter_enable :  STD_LOGIC;
                signal OpenMAC_0_CMP_arb_share_counter :  STD_LOGIC;
                signal OpenMAC_0_CMP_arb_share_counter_next_value :  STD_LOGIC;
                signal OpenMAC_0_CMP_arb_share_set_values :  STD_LOGIC;
                signal OpenMAC_0_CMP_beginbursttransfer_internal :  STD_LOGIC;
                signal OpenMAC_0_CMP_begins_xfer :  STD_LOGIC;
                signal OpenMAC_0_CMP_end_xfer :  STD_LOGIC;
                signal OpenMAC_0_CMP_firsttransfer :  STD_LOGIC;
                signal OpenMAC_0_CMP_grant_vector :  STD_LOGIC;
                signal OpenMAC_0_CMP_in_a_read_cycle :  STD_LOGIC;
                signal OpenMAC_0_CMP_in_a_write_cycle :  STD_LOGIC;
                signal OpenMAC_0_CMP_master_qreq_vector :  STD_LOGIC;
                signal OpenMAC_0_CMP_non_bursting_master_requests :  STD_LOGIC;
                signal OpenMAC_0_CMP_reg_firsttransfer :  STD_LOGIC;
                signal OpenMAC_0_CMP_slavearbiterlockenable :  STD_LOGIC;
                signal OpenMAC_0_CMP_slavearbiterlockenable2 :  STD_LOGIC;
                signal OpenMAC_0_CMP_unreg_firsttransfer :  STD_LOGIC;
                signal OpenMAC_0_CMP_waits_for_read :  STD_LOGIC;
                signal OpenMAC_0_CMP_waits_for_write :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_OpenMAC_0_CMP :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_niosII_openMac_clock_1_out_granted_OpenMAC_0_CMP :  STD_LOGIC;
                signal internal_niosII_openMac_clock_1_out_qualified_request_OpenMAC_0_CMP :  STD_LOGIC;
                signal internal_niosII_openMac_clock_1_out_requests_OpenMAC_0_CMP :  STD_LOGIC;
                signal niosII_openMac_clock_1_out_arbiterlock :  STD_LOGIC;
                signal niosII_openMac_clock_1_out_arbiterlock2 :  STD_LOGIC;
                signal niosII_openMac_clock_1_out_continuerequest :  STD_LOGIC;
                signal niosII_openMac_clock_1_out_saved_grant_OpenMAC_0_CMP :  STD_LOGIC;
                signal shifted_address_to_OpenMAC_0_CMP_from_niosII_openMac_clock_1_out :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal wait_for_OpenMAC_0_CMP_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT OpenMAC_0_CMP_end_xfer;
    end if;

  end process;

  OpenMAC_0_CMP_begins_xfer <= NOT d1_reasons_to_wait AND (internal_niosII_openMac_clock_1_out_qualified_request_OpenMAC_0_CMP);
  --assign OpenMAC_0_CMP_readdata_from_sa = OpenMAC_0_CMP_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  OpenMAC_0_CMP_readdata_from_sa <= OpenMAC_0_CMP_readdata;
  internal_niosII_openMac_clock_1_out_requests_OpenMAC_0_CMP <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((niosII_openMac_clock_1_out_read OR niosII_openMac_clock_1_out_write)))))));
  --OpenMAC_0_CMP_arb_share_counter set values, which is an e_mux
  OpenMAC_0_CMP_arb_share_set_values <= std_logic'('1');
  --OpenMAC_0_CMP_non_bursting_master_requests mux, which is an e_mux
  OpenMAC_0_CMP_non_bursting_master_requests <= internal_niosII_openMac_clock_1_out_requests_OpenMAC_0_CMP;
  --OpenMAC_0_CMP_any_bursting_master_saved_grant mux, which is an e_mux
  OpenMAC_0_CMP_any_bursting_master_saved_grant <= std_logic'('0');
  --OpenMAC_0_CMP_arb_share_counter_next_value assignment, which is an e_assign
  OpenMAC_0_CMP_arb_share_counter_next_value <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(OpenMAC_0_CMP_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(OpenMAC_0_CMP_arb_share_set_values))) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(OpenMAC_0_CMP_arb_share_counter) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(OpenMAC_0_CMP_arb_share_counter))) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))));
  --OpenMAC_0_CMP_allgrants all slave grants, which is an e_mux
  OpenMAC_0_CMP_allgrants <= OpenMAC_0_CMP_grant_vector;
  --OpenMAC_0_CMP_end_xfer assignment, which is an e_assign
  OpenMAC_0_CMP_end_xfer <= NOT ((OpenMAC_0_CMP_waits_for_read OR OpenMAC_0_CMP_waits_for_write));
  --end_xfer_arb_share_counter_term_OpenMAC_0_CMP arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_OpenMAC_0_CMP <= OpenMAC_0_CMP_end_xfer AND (((NOT OpenMAC_0_CMP_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --OpenMAC_0_CMP_arb_share_counter arbitration counter enable, which is an e_assign
  OpenMAC_0_CMP_arb_counter_enable <= ((end_xfer_arb_share_counter_term_OpenMAC_0_CMP AND OpenMAC_0_CMP_allgrants)) OR ((end_xfer_arb_share_counter_term_OpenMAC_0_CMP AND NOT OpenMAC_0_CMP_non_bursting_master_requests));
  --OpenMAC_0_CMP_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      OpenMAC_0_CMP_arb_share_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(OpenMAC_0_CMP_arb_counter_enable) = '1' then 
        OpenMAC_0_CMP_arb_share_counter <= OpenMAC_0_CMP_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --OpenMAC_0_CMP_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      OpenMAC_0_CMP_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((OpenMAC_0_CMP_master_qreq_vector AND end_xfer_arb_share_counter_term_OpenMAC_0_CMP)) OR ((end_xfer_arb_share_counter_term_OpenMAC_0_CMP AND NOT OpenMAC_0_CMP_non_bursting_master_requests)))) = '1' then 
        OpenMAC_0_CMP_slavearbiterlockenable <= OpenMAC_0_CMP_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --niosII_openMac_clock_1/out OpenMAC_0/CMP arbiterlock, which is an e_assign
  niosII_openMac_clock_1_out_arbiterlock <= OpenMAC_0_CMP_slavearbiterlockenable AND niosII_openMac_clock_1_out_continuerequest;
  --OpenMAC_0_CMP_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  OpenMAC_0_CMP_slavearbiterlockenable2 <= OpenMAC_0_CMP_arb_share_counter_next_value;
  --niosII_openMac_clock_1/out OpenMAC_0/CMP arbiterlock2, which is an e_assign
  niosII_openMac_clock_1_out_arbiterlock2 <= OpenMAC_0_CMP_slavearbiterlockenable2 AND niosII_openMac_clock_1_out_continuerequest;
  --OpenMAC_0_CMP_any_continuerequest at least one master continues requesting, which is an e_assign
  OpenMAC_0_CMP_any_continuerequest <= std_logic'('1');
  --niosII_openMac_clock_1_out_continuerequest continued request, which is an e_assign
  niosII_openMac_clock_1_out_continuerequest <= std_logic'('1');
  internal_niosII_openMac_clock_1_out_qualified_request_OpenMAC_0_CMP <= internal_niosII_openMac_clock_1_out_requests_OpenMAC_0_CMP;
  --OpenMAC_0_CMP_writedata mux, which is an e_mux
  OpenMAC_0_CMP_writedata <= niosII_openMac_clock_1_out_writedata;
  --master is always granted when requested
  internal_niosII_openMac_clock_1_out_granted_OpenMAC_0_CMP <= internal_niosII_openMac_clock_1_out_qualified_request_OpenMAC_0_CMP;
  --niosII_openMac_clock_1/out saved-grant OpenMAC_0/CMP, which is an e_assign
  niosII_openMac_clock_1_out_saved_grant_OpenMAC_0_CMP <= internal_niosII_openMac_clock_1_out_requests_OpenMAC_0_CMP;
  --allow new arb cycle for OpenMAC_0/CMP, which is an e_assign
  OpenMAC_0_CMP_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  OpenMAC_0_CMP_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  OpenMAC_0_CMP_master_qreq_vector <= std_logic'('1');
  --OpenMAC_0_CMP_reset_n assignment, which is an e_assign
  OpenMAC_0_CMP_reset_n <= reset_n;
  OpenMAC_0_CMP_chipselect <= internal_niosII_openMac_clock_1_out_granted_OpenMAC_0_CMP;
  --OpenMAC_0_CMP_firsttransfer first transaction, which is an e_assign
  OpenMAC_0_CMP_firsttransfer <= A_WE_StdLogic((std_logic'(OpenMAC_0_CMP_begins_xfer) = '1'), OpenMAC_0_CMP_unreg_firsttransfer, OpenMAC_0_CMP_reg_firsttransfer);
  --OpenMAC_0_CMP_unreg_firsttransfer first transaction, which is an e_assign
  OpenMAC_0_CMP_unreg_firsttransfer <= NOT ((OpenMAC_0_CMP_slavearbiterlockenable AND OpenMAC_0_CMP_any_continuerequest));
  --OpenMAC_0_CMP_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      OpenMAC_0_CMP_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(OpenMAC_0_CMP_begins_xfer) = '1' then 
        OpenMAC_0_CMP_reg_firsttransfer <= OpenMAC_0_CMP_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --OpenMAC_0_CMP_beginbursttransfer_internal begin burst transfer, which is an e_assign
  OpenMAC_0_CMP_beginbursttransfer_internal <= OpenMAC_0_CMP_begins_xfer;
  --~OpenMAC_0_CMP_read_n assignment, which is an e_mux
  OpenMAC_0_CMP_read_n <= NOT ((internal_niosII_openMac_clock_1_out_granted_OpenMAC_0_CMP AND niosII_openMac_clock_1_out_read));
  --~OpenMAC_0_CMP_write_n assignment, which is an e_mux
  OpenMAC_0_CMP_write_n <= NOT ((internal_niosII_openMac_clock_1_out_granted_OpenMAC_0_CMP AND niosII_openMac_clock_1_out_write));
  shifted_address_to_OpenMAC_0_CMP_from_niosII_openMac_clock_1_out <= niosII_openMac_clock_1_out_address_to_slave;
  --OpenMAC_0_CMP_address mux, which is an e_mux
  OpenMAC_0_CMP_address <= Vector_To_Std_Logic(A_SRL(shifted_address_to_OpenMAC_0_CMP_from_niosII_openMac_clock_1_out,std_logic_vector'("00000000000000000000000000000010")));
  --d1_OpenMAC_0_CMP_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_OpenMAC_0_CMP_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_OpenMAC_0_CMP_end_xfer <= OpenMAC_0_CMP_end_xfer;
    end if;

  end process;

  --OpenMAC_0_CMP_waits_for_read in a cycle, which is an e_mux
  OpenMAC_0_CMP_waits_for_read <= OpenMAC_0_CMP_in_a_read_cycle AND OpenMAC_0_CMP_begins_xfer;
  --OpenMAC_0_CMP_in_a_read_cycle assignment, which is an e_assign
  OpenMAC_0_CMP_in_a_read_cycle <= internal_niosII_openMac_clock_1_out_granted_OpenMAC_0_CMP AND niosII_openMac_clock_1_out_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= OpenMAC_0_CMP_in_a_read_cycle;
  --OpenMAC_0_CMP_waits_for_write in a cycle, which is an e_mux
  OpenMAC_0_CMP_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(OpenMAC_0_CMP_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --OpenMAC_0_CMP_in_a_write_cycle assignment, which is an e_assign
  OpenMAC_0_CMP_in_a_write_cycle <= internal_niosII_openMac_clock_1_out_granted_OpenMAC_0_CMP AND niosII_openMac_clock_1_out_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= OpenMAC_0_CMP_in_a_write_cycle;
  wait_for_OpenMAC_0_CMP_counter <= std_logic'('0');
  --~OpenMAC_0_CMP_byteenable_n byte enable port mux, which is an e_mux
  OpenMAC_0_CMP_byteenable_n <= A_EXT (NOT (A_WE_StdLogicVector((std_logic'((internal_niosII_openMac_clock_1_out_granted_OpenMAC_0_CMP)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (niosII_openMac_clock_1_out_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001")))), 4);
  --assign OpenMAC_0_CMP_irq_from_sa = OpenMAC_0_CMP_irq so that symbol knows where to group signals which may go to master only, which is an e_assign
  OpenMAC_0_CMP_irq_from_sa <= OpenMAC_0_CMP_irq;
  --vhdl renameroo for output signals
  niosII_openMac_clock_1_out_granted_OpenMAC_0_CMP <= internal_niosII_openMac_clock_1_out_granted_OpenMAC_0_CMP;
  --vhdl renameroo for output signals
  niosII_openMac_clock_1_out_qualified_request_OpenMAC_0_CMP <= internal_niosII_openMac_clock_1_out_qualified_request_OpenMAC_0_CMP;
  --vhdl renameroo for output signals
  niosII_openMac_clock_1_out_requests_OpenMAC_0_CMP <= internal_niosII_openMac_clock_1_out_requests_OpenMAC_0_CMP;
--synthesis translate_off
    --OpenMAC_0/CMP enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity OpenMAC_0_REG_arbitrator is 
        port (
              -- inputs:
                 signal OpenMAC_0_REG_irq : IN STD_LOGIC;
                 signal OpenMAC_0_REG_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal clk : IN STD_LOGIC;
                 signal niosII_openMac_clock_2_out_address_to_slave : IN STD_LOGIC_VECTOR (12 DOWNTO 0);
                 signal niosII_openMac_clock_2_out_byteenable : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal niosII_openMac_clock_2_out_read : IN STD_LOGIC;
                 signal niosII_openMac_clock_2_out_write : IN STD_LOGIC;
                 signal niosII_openMac_clock_2_out_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal OpenMAC_0_REG_address : OUT STD_LOGIC_VECTOR (11 DOWNTO 0);
                 signal OpenMAC_0_REG_byteenable_n : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal OpenMAC_0_REG_chipselect : OUT STD_LOGIC;
                 signal OpenMAC_0_REG_irq_from_sa : OUT STD_LOGIC;
                 signal OpenMAC_0_REG_read_n : OUT STD_LOGIC;
                 signal OpenMAC_0_REG_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal OpenMAC_0_REG_write_n : OUT STD_LOGIC;
                 signal OpenMAC_0_REG_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal d1_OpenMAC_0_REG_end_xfer : OUT STD_LOGIC;
                 signal niosII_openMac_clock_2_out_granted_OpenMAC_0_REG : OUT STD_LOGIC;
                 signal niosII_openMac_clock_2_out_qualified_request_OpenMAC_0_REG : OUT STD_LOGIC;
                 signal niosII_openMac_clock_2_out_read_data_valid_OpenMAC_0_REG : OUT STD_LOGIC;
                 signal niosII_openMac_clock_2_out_requests_OpenMAC_0_REG : OUT STD_LOGIC
              );
end entity OpenMAC_0_REG_arbitrator;


architecture europa of OpenMAC_0_REG_arbitrator is
                signal OpenMAC_0_REG_allgrants :  STD_LOGIC;
                signal OpenMAC_0_REG_allow_new_arb_cycle :  STD_LOGIC;
                signal OpenMAC_0_REG_any_bursting_master_saved_grant :  STD_LOGIC;
                signal OpenMAC_0_REG_any_continuerequest :  STD_LOGIC;
                signal OpenMAC_0_REG_arb_counter_enable :  STD_LOGIC;
                signal OpenMAC_0_REG_arb_share_counter :  STD_LOGIC;
                signal OpenMAC_0_REG_arb_share_counter_next_value :  STD_LOGIC;
                signal OpenMAC_0_REG_arb_share_set_values :  STD_LOGIC;
                signal OpenMAC_0_REG_beginbursttransfer_internal :  STD_LOGIC;
                signal OpenMAC_0_REG_begins_xfer :  STD_LOGIC;
                signal OpenMAC_0_REG_end_xfer :  STD_LOGIC;
                signal OpenMAC_0_REG_firsttransfer :  STD_LOGIC;
                signal OpenMAC_0_REG_grant_vector :  STD_LOGIC;
                signal OpenMAC_0_REG_in_a_read_cycle :  STD_LOGIC;
                signal OpenMAC_0_REG_in_a_write_cycle :  STD_LOGIC;
                signal OpenMAC_0_REG_master_qreq_vector :  STD_LOGIC;
                signal OpenMAC_0_REG_non_bursting_master_requests :  STD_LOGIC;
                signal OpenMAC_0_REG_reg_firsttransfer :  STD_LOGIC;
                signal OpenMAC_0_REG_slavearbiterlockenable :  STD_LOGIC;
                signal OpenMAC_0_REG_slavearbiterlockenable2 :  STD_LOGIC;
                signal OpenMAC_0_REG_unreg_firsttransfer :  STD_LOGIC;
                signal OpenMAC_0_REG_waits_for_read :  STD_LOGIC;
                signal OpenMAC_0_REG_waits_for_write :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_OpenMAC_0_REG :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_niosII_openMac_clock_2_out_granted_OpenMAC_0_REG :  STD_LOGIC;
                signal internal_niosII_openMac_clock_2_out_qualified_request_OpenMAC_0_REG :  STD_LOGIC;
                signal internal_niosII_openMac_clock_2_out_requests_OpenMAC_0_REG :  STD_LOGIC;
                signal niosII_openMac_clock_2_out_arbiterlock :  STD_LOGIC;
                signal niosII_openMac_clock_2_out_arbiterlock2 :  STD_LOGIC;
                signal niosII_openMac_clock_2_out_continuerequest :  STD_LOGIC;
                signal niosII_openMac_clock_2_out_saved_grant_OpenMAC_0_REG :  STD_LOGIC;
                signal shifted_address_to_OpenMAC_0_REG_from_niosII_openMac_clock_2_out :  STD_LOGIC_VECTOR (12 DOWNTO 0);
                signal wait_for_OpenMAC_0_REG_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT OpenMAC_0_REG_end_xfer;
    end if;

  end process;

  OpenMAC_0_REG_begins_xfer <= NOT d1_reasons_to_wait AND (internal_niosII_openMac_clock_2_out_qualified_request_OpenMAC_0_REG);
  --assign OpenMAC_0_REG_readdata_from_sa = OpenMAC_0_REG_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  OpenMAC_0_REG_readdata_from_sa <= OpenMAC_0_REG_readdata;
  internal_niosII_openMac_clock_2_out_requests_OpenMAC_0_REG <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((niosII_openMac_clock_2_out_read OR niosII_openMac_clock_2_out_write)))))));
  --OpenMAC_0_REG_arb_share_counter set values, which is an e_mux
  OpenMAC_0_REG_arb_share_set_values <= std_logic'('1');
  --OpenMAC_0_REG_non_bursting_master_requests mux, which is an e_mux
  OpenMAC_0_REG_non_bursting_master_requests <= internal_niosII_openMac_clock_2_out_requests_OpenMAC_0_REG;
  --OpenMAC_0_REG_any_bursting_master_saved_grant mux, which is an e_mux
  OpenMAC_0_REG_any_bursting_master_saved_grant <= std_logic'('0');
  --OpenMAC_0_REG_arb_share_counter_next_value assignment, which is an e_assign
  OpenMAC_0_REG_arb_share_counter_next_value <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(OpenMAC_0_REG_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(OpenMAC_0_REG_arb_share_set_values))) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(OpenMAC_0_REG_arb_share_counter) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(OpenMAC_0_REG_arb_share_counter))) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))));
  --OpenMAC_0_REG_allgrants all slave grants, which is an e_mux
  OpenMAC_0_REG_allgrants <= OpenMAC_0_REG_grant_vector;
  --OpenMAC_0_REG_end_xfer assignment, which is an e_assign
  OpenMAC_0_REG_end_xfer <= NOT ((OpenMAC_0_REG_waits_for_read OR OpenMAC_0_REG_waits_for_write));
  --end_xfer_arb_share_counter_term_OpenMAC_0_REG arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_OpenMAC_0_REG <= OpenMAC_0_REG_end_xfer AND (((NOT OpenMAC_0_REG_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --OpenMAC_0_REG_arb_share_counter arbitration counter enable, which is an e_assign
  OpenMAC_0_REG_arb_counter_enable <= ((end_xfer_arb_share_counter_term_OpenMAC_0_REG AND OpenMAC_0_REG_allgrants)) OR ((end_xfer_arb_share_counter_term_OpenMAC_0_REG AND NOT OpenMAC_0_REG_non_bursting_master_requests));
  --OpenMAC_0_REG_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      OpenMAC_0_REG_arb_share_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(OpenMAC_0_REG_arb_counter_enable) = '1' then 
        OpenMAC_0_REG_arb_share_counter <= OpenMAC_0_REG_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --OpenMAC_0_REG_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      OpenMAC_0_REG_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((OpenMAC_0_REG_master_qreq_vector AND end_xfer_arb_share_counter_term_OpenMAC_0_REG)) OR ((end_xfer_arb_share_counter_term_OpenMAC_0_REG AND NOT OpenMAC_0_REG_non_bursting_master_requests)))) = '1' then 
        OpenMAC_0_REG_slavearbiterlockenable <= OpenMAC_0_REG_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --niosII_openMac_clock_2/out OpenMAC_0/REG arbiterlock, which is an e_assign
  niosII_openMac_clock_2_out_arbiterlock <= OpenMAC_0_REG_slavearbiterlockenable AND niosII_openMac_clock_2_out_continuerequest;
  --OpenMAC_0_REG_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  OpenMAC_0_REG_slavearbiterlockenable2 <= OpenMAC_0_REG_arb_share_counter_next_value;
  --niosII_openMac_clock_2/out OpenMAC_0/REG arbiterlock2, which is an e_assign
  niosII_openMac_clock_2_out_arbiterlock2 <= OpenMAC_0_REG_slavearbiterlockenable2 AND niosII_openMac_clock_2_out_continuerequest;
  --OpenMAC_0_REG_any_continuerequest at least one master continues requesting, which is an e_assign
  OpenMAC_0_REG_any_continuerequest <= std_logic'('1');
  --niosII_openMac_clock_2_out_continuerequest continued request, which is an e_assign
  niosII_openMac_clock_2_out_continuerequest <= std_logic'('1');
  internal_niosII_openMac_clock_2_out_qualified_request_OpenMAC_0_REG <= internal_niosII_openMac_clock_2_out_requests_OpenMAC_0_REG;
  --OpenMAC_0_REG_writedata mux, which is an e_mux
  OpenMAC_0_REG_writedata <= niosII_openMac_clock_2_out_writedata;
  --master is always granted when requested
  internal_niosII_openMac_clock_2_out_granted_OpenMAC_0_REG <= internal_niosII_openMac_clock_2_out_qualified_request_OpenMAC_0_REG;
  --niosII_openMac_clock_2/out saved-grant OpenMAC_0/REG, which is an e_assign
  niosII_openMac_clock_2_out_saved_grant_OpenMAC_0_REG <= internal_niosII_openMac_clock_2_out_requests_OpenMAC_0_REG;
  --allow new arb cycle for OpenMAC_0/REG, which is an e_assign
  OpenMAC_0_REG_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  OpenMAC_0_REG_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  OpenMAC_0_REG_master_qreq_vector <= std_logic'('1');
  OpenMAC_0_REG_chipselect <= internal_niosII_openMac_clock_2_out_granted_OpenMAC_0_REG;
  --OpenMAC_0_REG_firsttransfer first transaction, which is an e_assign
  OpenMAC_0_REG_firsttransfer <= A_WE_StdLogic((std_logic'(OpenMAC_0_REG_begins_xfer) = '1'), OpenMAC_0_REG_unreg_firsttransfer, OpenMAC_0_REG_reg_firsttransfer);
  --OpenMAC_0_REG_unreg_firsttransfer first transaction, which is an e_assign
  OpenMAC_0_REG_unreg_firsttransfer <= NOT ((OpenMAC_0_REG_slavearbiterlockenable AND OpenMAC_0_REG_any_continuerequest));
  --OpenMAC_0_REG_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      OpenMAC_0_REG_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(OpenMAC_0_REG_begins_xfer) = '1' then 
        OpenMAC_0_REG_reg_firsttransfer <= OpenMAC_0_REG_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --OpenMAC_0_REG_beginbursttransfer_internal begin burst transfer, which is an e_assign
  OpenMAC_0_REG_beginbursttransfer_internal <= OpenMAC_0_REG_begins_xfer;
  --~OpenMAC_0_REG_read_n assignment, which is an e_mux
  OpenMAC_0_REG_read_n <= NOT ((internal_niosII_openMac_clock_2_out_granted_OpenMAC_0_REG AND niosII_openMac_clock_2_out_read));
  --~OpenMAC_0_REG_write_n assignment, which is an e_mux
  OpenMAC_0_REG_write_n <= NOT ((internal_niosII_openMac_clock_2_out_granted_OpenMAC_0_REG AND niosII_openMac_clock_2_out_write));
  shifted_address_to_OpenMAC_0_REG_from_niosII_openMac_clock_2_out <= niosII_openMac_clock_2_out_address_to_slave;
  --OpenMAC_0_REG_address mux, which is an e_mux
  OpenMAC_0_REG_address <= A_EXT (A_SRL(shifted_address_to_OpenMAC_0_REG_from_niosII_openMac_clock_2_out,std_logic_vector'("00000000000000000000000000000001")), 12);
  --d1_OpenMAC_0_REG_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_OpenMAC_0_REG_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_OpenMAC_0_REG_end_xfer <= OpenMAC_0_REG_end_xfer;
    end if;

  end process;

  --OpenMAC_0_REG_waits_for_read in a cycle, which is an e_mux
  OpenMAC_0_REG_waits_for_read <= OpenMAC_0_REG_in_a_read_cycle AND OpenMAC_0_REG_begins_xfer;
  --OpenMAC_0_REG_in_a_read_cycle assignment, which is an e_assign
  OpenMAC_0_REG_in_a_read_cycle <= internal_niosII_openMac_clock_2_out_granted_OpenMAC_0_REG AND niosII_openMac_clock_2_out_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= OpenMAC_0_REG_in_a_read_cycle;
  --OpenMAC_0_REG_waits_for_write in a cycle, which is an e_mux
  OpenMAC_0_REG_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(OpenMAC_0_REG_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --OpenMAC_0_REG_in_a_write_cycle assignment, which is an e_assign
  OpenMAC_0_REG_in_a_write_cycle <= internal_niosII_openMac_clock_2_out_granted_OpenMAC_0_REG AND niosII_openMac_clock_2_out_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= OpenMAC_0_REG_in_a_write_cycle;
  wait_for_OpenMAC_0_REG_counter <= std_logic'('0');
  --~OpenMAC_0_REG_byteenable_n byte enable port mux, which is an e_mux
  OpenMAC_0_REG_byteenable_n <= A_EXT (NOT (A_WE_StdLogicVector((std_logic'((internal_niosII_openMac_clock_2_out_granted_OpenMAC_0_REG)) = '1'), (std_logic_vector'("000000000000000000000000000000") & (niosII_openMac_clock_2_out_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001")))), 2);
  --assign OpenMAC_0_REG_irq_from_sa = OpenMAC_0_REG_irq so that symbol knows where to group signals which may go to master only, which is an e_assign
  OpenMAC_0_REG_irq_from_sa <= OpenMAC_0_REG_irq;
  --vhdl renameroo for output signals
  niosII_openMac_clock_2_out_granted_OpenMAC_0_REG <= internal_niosII_openMac_clock_2_out_granted_OpenMAC_0_REG;
  --vhdl renameroo for output signals
  niosII_openMac_clock_2_out_qualified_request_OpenMAC_0_REG <= internal_niosII_openMac_clock_2_out_qualified_request_OpenMAC_0_REG;
  --vhdl renameroo for output signals
  niosII_openMac_clock_2_out_requests_OpenMAC_0_REG <= internal_niosII_openMac_clock_2_out_requests_OpenMAC_0_REG;
--synthesis translate_off
    --OpenMAC_0/REG enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity OpenMAC_0_iBuf_arbitrator is 
        port (
              -- inputs:
                 signal OpenMAC_0_iBuf_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal clk : IN STD_LOGIC;
                 signal pcp_cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (25 DOWNTO 0);
                 signal pcp_cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal pcp_cpu_data_master_read : IN STD_LOGIC;
                 signal pcp_cpu_data_master_waitrequest : IN STD_LOGIC;
                 signal pcp_cpu_data_master_write : IN STD_LOGIC;
                 signal pcp_cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal OpenMAC_0_iBuf_address : OUT STD_LOGIC_VECTOR (12 DOWNTO 0);
                 signal OpenMAC_0_iBuf_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal OpenMAC_0_iBuf_chipselect : OUT STD_LOGIC;
                 signal OpenMAC_0_iBuf_read_n : OUT STD_LOGIC;
                 signal OpenMAC_0_iBuf_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal OpenMAC_0_iBuf_wait_counter_eq_0 : OUT STD_LOGIC;
                 signal OpenMAC_0_iBuf_write_n : OUT STD_LOGIC;
                 signal OpenMAC_0_iBuf_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal d1_OpenMAC_0_iBuf_end_xfer : OUT STD_LOGIC;
                 signal pcp_cpu_data_master_granted_OpenMAC_0_iBuf : OUT STD_LOGIC;
                 signal pcp_cpu_data_master_qualified_request_OpenMAC_0_iBuf : OUT STD_LOGIC;
                 signal pcp_cpu_data_master_read_data_valid_OpenMAC_0_iBuf : OUT STD_LOGIC;
                 signal pcp_cpu_data_master_requests_OpenMAC_0_iBuf : OUT STD_LOGIC
              );
end entity OpenMAC_0_iBuf_arbitrator;


architecture europa of OpenMAC_0_iBuf_arbitrator is
                signal OpenMAC_0_iBuf_allgrants :  STD_LOGIC;
                signal OpenMAC_0_iBuf_allow_new_arb_cycle :  STD_LOGIC;
                signal OpenMAC_0_iBuf_any_bursting_master_saved_grant :  STD_LOGIC;
                signal OpenMAC_0_iBuf_any_continuerequest :  STD_LOGIC;
                signal OpenMAC_0_iBuf_arb_counter_enable :  STD_LOGIC;
                signal OpenMAC_0_iBuf_arb_share_counter :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal OpenMAC_0_iBuf_arb_share_counter_next_value :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal OpenMAC_0_iBuf_arb_share_set_values :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal OpenMAC_0_iBuf_beginbursttransfer_internal :  STD_LOGIC;
                signal OpenMAC_0_iBuf_begins_xfer :  STD_LOGIC;
                signal OpenMAC_0_iBuf_counter_load_value :  STD_LOGIC;
                signal OpenMAC_0_iBuf_end_xfer :  STD_LOGIC;
                signal OpenMAC_0_iBuf_firsttransfer :  STD_LOGIC;
                signal OpenMAC_0_iBuf_grant_vector :  STD_LOGIC;
                signal OpenMAC_0_iBuf_in_a_read_cycle :  STD_LOGIC;
                signal OpenMAC_0_iBuf_in_a_write_cycle :  STD_LOGIC;
                signal OpenMAC_0_iBuf_master_qreq_vector :  STD_LOGIC;
                signal OpenMAC_0_iBuf_non_bursting_master_requests :  STD_LOGIC;
                signal OpenMAC_0_iBuf_reg_firsttransfer :  STD_LOGIC;
                signal OpenMAC_0_iBuf_slavearbiterlockenable :  STD_LOGIC;
                signal OpenMAC_0_iBuf_slavearbiterlockenable2 :  STD_LOGIC;
                signal OpenMAC_0_iBuf_unreg_firsttransfer :  STD_LOGIC;
                signal OpenMAC_0_iBuf_wait_counter :  STD_LOGIC;
                signal OpenMAC_0_iBuf_waits_for_read :  STD_LOGIC;
                signal OpenMAC_0_iBuf_waits_for_write :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_OpenMAC_0_iBuf :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_OpenMAC_0_iBuf_wait_counter_eq_0 :  STD_LOGIC;
                signal internal_pcp_cpu_data_master_granted_OpenMAC_0_iBuf :  STD_LOGIC;
                signal internal_pcp_cpu_data_master_qualified_request_OpenMAC_0_iBuf :  STD_LOGIC;
                signal internal_pcp_cpu_data_master_requests_OpenMAC_0_iBuf :  STD_LOGIC;
                signal pcp_cpu_data_master_arbiterlock :  STD_LOGIC;
                signal pcp_cpu_data_master_arbiterlock2 :  STD_LOGIC;
                signal pcp_cpu_data_master_continuerequest :  STD_LOGIC;
                signal pcp_cpu_data_master_saved_grant_OpenMAC_0_iBuf :  STD_LOGIC;
                signal shifted_address_to_OpenMAC_0_iBuf_from_pcp_cpu_data_master :  STD_LOGIC_VECTOR (25 DOWNTO 0);
                signal wait_for_OpenMAC_0_iBuf_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT OpenMAC_0_iBuf_end_xfer;
    end if;

  end process;

  OpenMAC_0_iBuf_begins_xfer <= NOT d1_reasons_to_wait AND (internal_pcp_cpu_data_master_qualified_request_OpenMAC_0_iBuf);
  --assign OpenMAC_0_iBuf_readdata_from_sa = OpenMAC_0_iBuf_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  OpenMAC_0_iBuf_readdata_from_sa <= OpenMAC_0_iBuf_readdata;
  internal_pcp_cpu_data_master_requests_OpenMAC_0_iBuf <= to_std_logic(((Std_Logic_Vector'(pcp_cpu_data_master_address_to_slave(25 DOWNTO 15) & std_logic_vector'("000000000000000")) = std_logic_vector'("00000000001000000000000000")))) AND ((pcp_cpu_data_master_read OR pcp_cpu_data_master_write));
  --OpenMAC_0_iBuf_arb_share_counter set values, which is an e_mux
  OpenMAC_0_iBuf_arb_share_set_values <= std_logic_vector'("01");
  --OpenMAC_0_iBuf_non_bursting_master_requests mux, which is an e_mux
  OpenMAC_0_iBuf_non_bursting_master_requests <= internal_pcp_cpu_data_master_requests_OpenMAC_0_iBuf;
  --OpenMAC_0_iBuf_any_bursting_master_saved_grant mux, which is an e_mux
  OpenMAC_0_iBuf_any_bursting_master_saved_grant <= std_logic'('0');
  --OpenMAC_0_iBuf_arb_share_counter_next_value assignment, which is an e_assign
  OpenMAC_0_iBuf_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(OpenMAC_0_iBuf_firsttransfer) = '1'), (((std_logic_vector'("0000000000000000000000000000000") & (OpenMAC_0_iBuf_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(OpenMAC_0_iBuf_arb_share_counter)) = '1'), (((std_logic_vector'("0000000000000000000000000000000") & (OpenMAC_0_iBuf_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 2);
  --OpenMAC_0_iBuf_allgrants all slave grants, which is an e_mux
  OpenMAC_0_iBuf_allgrants <= OpenMAC_0_iBuf_grant_vector;
  --OpenMAC_0_iBuf_end_xfer assignment, which is an e_assign
  OpenMAC_0_iBuf_end_xfer <= NOT ((OpenMAC_0_iBuf_waits_for_read OR OpenMAC_0_iBuf_waits_for_write));
  --end_xfer_arb_share_counter_term_OpenMAC_0_iBuf arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_OpenMAC_0_iBuf <= OpenMAC_0_iBuf_end_xfer AND (((NOT OpenMAC_0_iBuf_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --OpenMAC_0_iBuf_arb_share_counter arbitration counter enable, which is an e_assign
  OpenMAC_0_iBuf_arb_counter_enable <= ((end_xfer_arb_share_counter_term_OpenMAC_0_iBuf AND OpenMAC_0_iBuf_allgrants)) OR ((end_xfer_arb_share_counter_term_OpenMAC_0_iBuf AND NOT OpenMAC_0_iBuf_non_bursting_master_requests));
  --OpenMAC_0_iBuf_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      OpenMAC_0_iBuf_arb_share_counter <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      if std_logic'(OpenMAC_0_iBuf_arb_counter_enable) = '1' then 
        OpenMAC_0_iBuf_arb_share_counter <= OpenMAC_0_iBuf_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --OpenMAC_0_iBuf_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      OpenMAC_0_iBuf_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((OpenMAC_0_iBuf_master_qreq_vector AND end_xfer_arb_share_counter_term_OpenMAC_0_iBuf)) OR ((end_xfer_arb_share_counter_term_OpenMAC_0_iBuf AND NOT OpenMAC_0_iBuf_non_bursting_master_requests)))) = '1' then 
        OpenMAC_0_iBuf_slavearbiterlockenable <= or_reduce(OpenMAC_0_iBuf_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --pcp_cpu/data_master OpenMAC_0/iBuf arbiterlock, which is an e_assign
  pcp_cpu_data_master_arbiterlock <= OpenMAC_0_iBuf_slavearbiterlockenable AND pcp_cpu_data_master_continuerequest;
  --OpenMAC_0_iBuf_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  OpenMAC_0_iBuf_slavearbiterlockenable2 <= or_reduce(OpenMAC_0_iBuf_arb_share_counter_next_value);
  --pcp_cpu/data_master OpenMAC_0/iBuf arbiterlock2, which is an e_assign
  pcp_cpu_data_master_arbiterlock2 <= OpenMAC_0_iBuf_slavearbiterlockenable2 AND pcp_cpu_data_master_continuerequest;
  --OpenMAC_0_iBuf_any_continuerequest at least one master continues requesting, which is an e_assign
  OpenMAC_0_iBuf_any_continuerequest <= std_logic'('1');
  --pcp_cpu_data_master_continuerequest continued request, which is an e_assign
  pcp_cpu_data_master_continuerequest <= std_logic'('1');
  internal_pcp_cpu_data_master_qualified_request_OpenMAC_0_iBuf <= internal_pcp_cpu_data_master_requests_OpenMAC_0_iBuf AND NOT (((NOT pcp_cpu_data_master_waitrequest) AND pcp_cpu_data_master_write));
  --OpenMAC_0_iBuf_writedata mux, which is an e_mux
  OpenMAC_0_iBuf_writedata <= pcp_cpu_data_master_writedata;
  --master is always granted when requested
  internal_pcp_cpu_data_master_granted_OpenMAC_0_iBuf <= internal_pcp_cpu_data_master_qualified_request_OpenMAC_0_iBuf;
  --pcp_cpu/data_master saved-grant OpenMAC_0/iBuf, which is an e_assign
  pcp_cpu_data_master_saved_grant_OpenMAC_0_iBuf <= internal_pcp_cpu_data_master_requests_OpenMAC_0_iBuf;
  --allow new arb cycle for OpenMAC_0/iBuf, which is an e_assign
  OpenMAC_0_iBuf_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  OpenMAC_0_iBuf_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  OpenMAC_0_iBuf_master_qreq_vector <= std_logic'('1');
  OpenMAC_0_iBuf_chipselect <= internal_pcp_cpu_data_master_granted_OpenMAC_0_iBuf;
  --OpenMAC_0_iBuf_firsttransfer first transaction, which is an e_assign
  OpenMAC_0_iBuf_firsttransfer <= A_WE_StdLogic((std_logic'(OpenMAC_0_iBuf_begins_xfer) = '1'), OpenMAC_0_iBuf_unreg_firsttransfer, OpenMAC_0_iBuf_reg_firsttransfer);
  --OpenMAC_0_iBuf_unreg_firsttransfer first transaction, which is an e_assign
  OpenMAC_0_iBuf_unreg_firsttransfer <= NOT ((OpenMAC_0_iBuf_slavearbiterlockenable AND OpenMAC_0_iBuf_any_continuerequest));
  --OpenMAC_0_iBuf_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      OpenMAC_0_iBuf_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(OpenMAC_0_iBuf_begins_xfer) = '1' then 
        OpenMAC_0_iBuf_reg_firsttransfer <= OpenMAC_0_iBuf_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --OpenMAC_0_iBuf_beginbursttransfer_internal begin burst transfer, which is an e_assign
  OpenMAC_0_iBuf_beginbursttransfer_internal <= OpenMAC_0_iBuf_begins_xfer;
  --~OpenMAC_0_iBuf_read_n assignment, which is an e_mux
  OpenMAC_0_iBuf_read_n <= NOT ((internal_pcp_cpu_data_master_granted_OpenMAC_0_iBuf AND pcp_cpu_data_master_read));
  --~OpenMAC_0_iBuf_write_n assignment, which is an e_mux
  OpenMAC_0_iBuf_write_n <= NOT ((internal_pcp_cpu_data_master_granted_OpenMAC_0_iBuf AND pcp_cpu_data_master_write));
  shifted_address_to_OpenMAC_0_iBuf_from_pcp_cpu_data_master <= pcp_cpu_data_master_address_to_slave;
  --OpenMAC_0_iBuf_address mux, which is an e_mux
  OpenMAC_0_iBuf_address <= A_EXT (A_SRL(shifted_address_to_OpenMAC_0_iBuf_from_pcp_cpu_data_master,std_logic_vector'("00000000000000000000000000000010")), 13);
  --d1_OpenMAC_0_iBuf_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_OpenMAC_0_iBuf_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_OpenMAC_0_iBuf_end_xfer <= OpenMAC_0_iBuf_end_xfer;
    end if;

  end process;

  --OpenMAC_0_iBuf_waits_for_read in a cycle, which is an e_mux
  OpenMAC_0_iBuf_waits_for_read <= OpenMAC_0_iBuf_in_a_read_cycle AND wait_for_OpenMAC_0_iBuf_counter;
  --OpenMAC_0_iBuf_in_a_read_cycle assignment, which is an e_assign
  OpenMAC_0_iBuf_in_a_read_cycle <= internal_pcp_cpu_data_master_granted_OpenMAC_0_iBuf AND pcp_cpu_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= OpenMAC_0_iBuf_in_a_read_cycle;
  --OpenMAC_0_iBuf_waits_for_write in a cycle, which is an e_mux
  OpenMAC_0_iBuf_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(OpenMAC_0_iBuf_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --OpenMAC_0_iBuf_in_a_write_cycle assignment, which is an e_assign
  OpenMAC_0_iBuf_in_a_write_cycle <= internal_pcp_cpu_data_master_granted_OpenMAC_0_iBuf AND pcp_cpu_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= OpenMAC_0_iBuf_in_a_write_cycle;
  internal_OpenMAC_0_iBuf_wait_counter_eq_0 <= to_std_logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(OpenMAC_0_iBuf_wait_counter))) = std_logic_vector'("00000000000000000000000000000000")));
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      OpenMAC_0_iBuf_wait_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      OpenMAC_0_iBuf_wait_counter <= OpenMAC_0_iBuf_counter_load_value;
    end if;

  end process;

  OpenMAC_0_iBuf_counter_load_value <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(((OpenMAC_0_iBuf_in_a_read_cycle AND OpenMAC_0_iBuf_begins_xfer))) = '1'), std_logic_vector'("000000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'((NOT internal_OpenMAC_0_iBuf_wait_counter_eq_0)) = '1'), ((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(OpenMAC_0_iBuf_wait_counter))) - std_logic_vector'("000000000000000000000000000000001")), std_logic_vector'("000000000000000000000000000000000"))));
  wait_for_OpenMAC_0_iBuf_counter <= OpenMAC_0_iBuf_begins_xfer OR NOT internal_OpenMAC_0_iBuf_wait_counter_eq_0;
  --OpenMAC_0_iBuf_byteenable byte enable port mux, which is an e_mux
  OpenMAC_0_iBuf_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_pcp_cpu_data_master_granted_OpenMAC_0_iBuf)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (pcp_cpu_data_master_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))), 4);
  --vhdl renameroo for output signals
  OpenMAC_0_iBuf_wait_counter_eq_0 <= internal_OpenMAC_0_iBuf_wait_counter_eq_0;
  --vhdl renameroo for output signals
  pcp_cpu_data_master_granted_OpenMAC_0_iBuf <= internal_pcp_cpu_data_master_granted_OpenMAC_0_iBuf;
  --vhdl renameroo for output signals
  pcp_cpu_data_master_qualified_request_OpenMAC_0_iBuf <= internal_pcp_cpu_data_master_qualified_request_OpenMAC_0_iBuf;
  --vhdl renameroo for output signals
  pcp_cpu_data_master_requests_OpenMAC_0_iBuf <= internal_pcp_cpu_data_master_requests_OpenMAC_0_iBuf;
--synthesis translate_off
    --OpenMAC_0/iBuf enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity altpll_0_pll_slave_arbitrator is 
        port (
              -- inputs:
                 signal altpll_0_pll_slave_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal clk : IN STD_LOGIC;
                 signal niosII_openMac_clock_3_out_address_to_slave : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal niosII_openMac_clock_3_out_read : IN STD_LOGIC;
                 signal niosII_openMac_clock_3_out_write : IN STD_LOGIC;
                 signal niosII_openMac_clock_3_out_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal altpll_0_pll_slave_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal altpll_0_pll_slave_read : OUT STD_LOGIC;
                 signal altpll_0_pll_slave_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal altpll_0_pll_slave_reset : OUT STD_LOGIC;
                 signal altpll_0_pll_slave_write : OUT STD_LOGIC;
                 signal altpll_0_pll_slave_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal d1_altpll_0_pll_slave_end_xfer : OUT STD_LOGIC;
                 signal niosII_openMac_clock_3_out_granted_altpll_0_pll_slave : OUT STD_LOGIC;
                 signal niosII_openMac_clock_3_out_qualified_request_altpll_0_pll_slave : OUT STD_LOGIC;
                 signal niosII_openMac_clock_3_out_read_data_valid_altpll_0_pll_slave : OUT STD_LOGIC;
                 signal niosII_openMac_clock_3_out_requests_altpll_0_pll_slave : OUT STD_LOGIC
              );
end entity altpll_0_pll_slave_arbitrator;


architecture europa of altpll_0_pll_slave_arbitrator is
                signal altpll_0_pll_slave_allgrants :  STD_LOGIC;
                signal altpll_0_pll_slave_allow_new_arb_cycle :  STD_LOGIC;
                signal altpll_0_pll_slave_any_bursting_master_saved_grant :  STD_LOGIC;
                signal altpll_0_pll_slave_any_continuerequest :  STD_LOGIC;
                signal altpll_0_pll_slave_arb_counter_enable :  STD_LOGIC;
                signal altpll_0_pll_slave_arb_share_counter :  STD_LOGIC;
                signal altpll_0_pll_slave_arb_share_counter_next_value :  STD_LOGIC;
                signal altpll_0_pll_slave_arb_share_set_values :  STD_LOGIC;
                signal altpll_0_pll_slave_beginbursttransfer_internal :  STD_LOGIC;
                signal altpll_0_pll_slave_begins_xfer :  STD_LOGIC;
                signal altpll_0_pll_slave_end_xfer :  STD_LOGIC;
                signal altpll_0_pll_slave_firsttransfer :  STD_LOGIC;
                signal altpll_0_pll_slave_grant_vector :  STD_LOGIC;
                signal altpll_0_pll_slave_in_a_read_cycle :  STD_LOGIC;
                signal altpll_0_pll_slave_in_a_write_cycle :  STD_LOGIC;
                signal altpll_0_pll_slave_master_qreq_vector :  STD_LOGIC;
                signal altpll_0_pll_slave_non_bursting_master_requests :  STD_LOGIC;
                signal altpll_0_pll_slave_reg_firsttransfer :  STD_LOGIC;
                signal altpll_0_pll_slave_slavearbiterlockenable :  STD_LOGIC;
                signal altpll_0_pll_slave_slavearbiterlockenable2 :  STD_LOGIC;
                signal altpll_0_pll_slave_unreg_firsttransfer :  STD_LOGIC;
                signal altpll_0_pll_slave_waits_for_read :  STD_LOGIC;
                signal altpll_0_pll_slave_waits_for_write :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_altpll_0_pll_slave :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_niosII_openMac_clock_3_out_granted_altpll_0_pll_slave :  STD_LOGIC;
                signal internal_niosII_openMac_clock_3_out_qualified_request_altpll_0_pll_slave :  STD_LOGIC;
                signal internal_niosII_openMac_clock_3_out_requests_altpll_0_pll_slave :  STD_LOGIC;
                signal niosII_openMac_clock_3_out_arbiterlock :  STD_LOGIC;
                signal niosII_openMac_clock_3_out_arbiterlock2 :  STD_LOGIC;
                signal niosII_openMac_clock_3_out_continuerequest :  STD_LOGIC;
                signal niosII_openMac_clock_3_out_saved_grant_altpll_0_pll_slave :  STD_LOGIC;
                signal shifted_address_to_altpll_0_pll_slave_from_niosII_openMac_clock_3_out :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal wait_for_altpll_0_pll_slave_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT altpll_0_pll_slave_end_xfer;
    end if;

  end process;

  altpll_0_pll_slave_begins_xfer <= NOT d1_reasons_to_wait AND (internal_niosII_openMac_clock_3_out_qualified_request_altpll_0_pll_slave);
  --assign altpll_0_pll_slave_readdata_from_sa = altpll_0_pll_slave_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  altpll_0_pll_slave_readdata_from_sa <= altpll_0_pll_slave_readdata;
  internal_niosII_openMac_clock_3_out_requests_altpll_0_pll_slave <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((niosII_openMac_clock_3_out_read OR niosII_openMac_clock_3_out_write)))))));
  --altpll_0_pll_slave_arb_share_counter set values, which is an e_mux
  altpll_0_pll_slave_arb_share_set_values <= std_logic'('1');
  --altpll_0_pll_slave_non_bursting_master_requests mux, which is an e_mux
  altpll_0_pll_slave_non_bursting_master_requests <= internal_niosII_openMac_clock_3_out_requests_altpll_0_pll_slave;
  --altpll_0_pll_slave_any_bursting_master_saved_grant mux, which is an e_mux
  altpll_0_pll_slave_any_bursting_master_saved_grant <= std_logic'('0');
  --altpll_0_pll_slave_arb_share_counter_next_value assignment, which is an e_assign
  altpll_0_pll_slave_arb_share_counter_next_value <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(altpll_0_pll_slave_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(altpll_0_pll_slave_arb_share_set_values))) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(altpll_0_pll_slave_arb_share_counter) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(altpll_0_pll_slave_arb_share_counter))) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))));
  --altpll_0_pll_slave_allgrants all slave grants, which is an e_mux
  altpll_0_pll_slave_allgrants <= altpll_0_pll_slave_grant_vector;
  --altpll_0_pll_slave_end_xfer assignment, which is an e_assign
  altpll_0_pll_slave_end_xfer <= NOT ((altpll_0_pll_slave_waits_for_read OR altpll_0_pll_slave_waits_for_write));
  --end_xfer_arb_share_counter_term_altpll_0_pll_slave arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_altpll_0_pll_slave <= altpll_0_pll_slave_end_xfer AND (((NOT altpll_0_pll_slave_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --altpll_0_pll_slave_arb_share_counter arbitration counter enable, which is an e_assign
  altpll_0_pll_slave_arb_counter_enable <= ((end_xfer_arb_share_counter_term_altpll_0_pll_slave AND altpll_0_pll_slave_allgrants)) OR ((end_xfer_arb_share_counter_term_altpll_0_pll_slave AND NOT altpll_0_pll_slave_non_bursting_master_requests));
  --altpll_0_pll_slave_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      altpll_0_pll_slave_arb_share_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(altpll_0_pll_slave_arb_counter_enable) = '1' then 
        altpll_0_pll_slave_arb_share_counter <= altpll_0_pll_slave_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --altpll_0_pll_slave_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      altpll_0_pll_slave_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((altpll_0_pll_slave_master_qreq_vector AND end_xfer_arb_share_counter_term_altpll_0_pll_slave)) OR ((end_xfer_arb_share_counter_term_altpll_0_pll_slave AND NOT altpll_0_pll_slave_non_bursting_master_requests)))) = '1' then 
        altpll_0_pll_slave_slavearbiterlockenable <= altpll_0_pll_slave_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --niosII_openMac_clock_3/out altpll_0/pll_slave arbiterlock, which is an e_assign
  niosII_openMac_clock_3_out_arbiterlock <= altpll_0_pll_slave_slavearbiterlockenable AND niosII_openMac_clock_3_out_continuerequest;
  --altpll_0_pll_slave_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  altpll_0_pll_slave_slavearbiterlockenable2 <= altpll_0_pll_slave_arb_share_counter_next_value;
  --niosII_openMac_clock_3/out altpll_0/pll_slave arbiterlock2, which is an e_assign
  niosII_openMac_clock_3_out_arbiterlock2 <= altpll_0_pll_slave_slavearbiterlockenable2 AND niosII_openMac_clock_3_out_continuerequest;
  --altpll_0_pll_slave_any_continuerequest at least one master continues requesting, which is an e_assign
  altpll_0_pll_slave_any_continuerequest <= std_logic'('1');
  --niosII_openMac_clock_3_out_continuerequest continued request, which is an e_assign
  niosII_openMac_clock_3_out_continuerequest <= std_logic'('1');
  internal_niosII_openMac_clock_3_out_qualified_request_altpll_0_pll_slave <= internal_niosII_openMac_clock_3_out_requests_altpll_0_pll_slave;
  --altpll_0_pll_slave_writedata mux, which is an e_mux
  altpll_0_pll_slave_writedata <= niosII_openMac_clock_3_out_writedata;
  --master is always granted when requested
  internal_niosII_openMac_clock_3_out_granted_altpll_0_pll_slave <= internal_niosII_openMac_clock_3_out_qualified_request_altpll_0_pll_slave;
  --niosII_openMac_clock_3/out saved-grant altpll_0/pll_slave, which is an e_assign
  niosII_openMac_clock_3_out_saved_grant_altpll_0_pll_slave <= internal_niosII_openMac_clock_3_out_requests_altpll_0_pll_slave;
  --allow new arb cycle for altpll_0/pll_slave, which is an e_assign
  altpll_0_pll_slave_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  altpll_0_pll_slave_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  altpll_0_pll_slave_master_qreq_vector <= std_logic'('1');
  --~altpll_0_pll_slave_reset assignment, which is an e_assign
  altpll_0_pll_slave_reset <= NOT reset_n;
  --altpll_0_pll_slave_firsttransfer first transaction, which is an e_assign
  altpll_0_pll_slave_firsttransfer <= A_WE_StdLogic((std_logic'(altpll_0_pll_slave_begins_xfer) = '1'), altpll_0_pll_slave_unreg_firsttransfer, altpll_0_pll_slave_reg_firsttransfer);
  --altpll_0_pll_slave_unreg_firsttransfer first transaction, which is an e_assign
  altpll_0_pll_slave_unreg_firsttransfer <= NOT ((altpll_0_pll_slave_slavearbiterlockenable AND altpll_0_pll_slave_any_continuerequest));
  --altpll_0_pll_slave_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      altpll_0_pll_slave_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(altpll_0_pll_slave_begins_xfer) = '1' then 
        altpll_0_pll_slave_reg_firsttransfer <= altpll_0_pll_slave_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --altpll_0_pll_slave_beginbursttransfer_internal begin burst transfer, which is an e_assign
  altpll_0_pll_slave_beginbursttransfer_internal <= altpll_0_pll_slave_begins_xfer;
  --altpll_0_pll_slave_read assignment, which is an e_mux
  altpll_0_pll_slave_read <= internal_niosII_openMac_clock_3_out_granted_altpll_0_pll_slave AND niosII_openMac_clock_3_out_read;
  --altpll_0_pll_slave_write assignment, which is an e_mux
  altpll_0_pll_slave_write <= internal_niosII_openMac_clock_3_out_granted_altpll_0_pll_slave AND niosII_openMac_clock_3_out_write;
  shifted_address_to_altpll_0_pll_slave_from_niosII_openMac_clock_3_out <= niosII_openMac_clock_3_out_address_to_slave;
  --altpll_0_pll_slave_address mux, which is an e_mux
  altpll_0_pll_slave_address <= A_EXT (A_SRL(shifted_address_to_altpll_0_pll_slave_from_niosII_openMac_clock_3_out,std_logic_vector'("00000000000000000000000000000010")), 2);
  --d1_altpll_0_pll_slave_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_altpll_0_pll_slave_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_altpll_0_pll_slave_end_xfer <= altpll_0_pll_slave_end_xfer;
    end if;

  end process;

  --altpll_0_pll_slave_waits_for_read in a cycle, which is an e_mux
  altpll_0_pll_slave_waits_for_read <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(altpll_0_pll_slave_in_a_read_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --altpll_0_pll_slave_in_a_read_cycle assignment, which is an e_assign
  altpll_0_pll_slave_in_a_read_cycle <= internal_niosII_openMac_clock_3_out_granted_altpll_0_pll_slave AND niosII_openMac_clock_3_out_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= altpll_0_pll_slave_in_a_read_cycle;
  --altpll_0_pll_slave_waits_for_write in a cycle, which is an e_mux
  altpll_0_pll_slave_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(altpll_0_pll_slave_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --altpll_0_pll_slave_in_a_write_cycle assignment, which is an e_assign
  altpll_0_pll_slave_in_a_write_cycle <= internal_niosII_openMac_clock_3_out_granted_altpll_0_pll_slave AND niosII_openMac_clock_3_out_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= altpll_0_pll_slave_in_a_write_cycle;
  wait_for_altpll_0_pll_slave_counter <= std_logic'('0');
  --vhdl renameroo for output signals
  niosII_openMac_clock_3_out_granted_altpll_0_pll_slave <= internal_niosII_openMac_clock_3_out_granted_altpll_0_pll_slave;
  --vhdl renameroo for output signals
  niosII_openMac_clock_3_out_qualified_request_altpll_0_pll_slave <= internal_niosII_openMac_clock_3_out_qualified_request_altpll_0_pll_slave;
  --vhdl renameroo for output signals
  niosII_openMac_clock_3_out_requests_altpll_0_pll_slave <= internal_niosII_openMac_clock_3_out_requests_altpll_0_pll_slave;
--synthesis translate_off
    --altpll_0/pll_slave enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity ap_cpu_jtag_debug_module_arbitrator is 
        port (
              -- inputs:
                 signal ap_cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (25 DOWNTO 0);
                 signal ap_cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal ap_cpu_data_master_debugaccess : IN STD_LOGIC;
                 signal ap_cpu_data_master_read : IN STD_LOGIC;
                 signal ap_cpu_data_master_waitrequest : IN STD_LOGIC;
                 signal ap_cpu_data_master_write : IN STD_LOGIC;
                 signal ap_cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal ap_cpu_instruction_master_address_to_slave : IN STD_LOGIC_VECTOR (25 DOWNTO 0);
                 signal ap_cpu_instruction_master_latency_counter : IN STD_LOGIC;
                 signal ap_cpu_instruction_master_read : IN STD_LOGIC;
                 signal ap_cpu_instruction_master_read_data_valid_sdram_0_s1_shift_register : IN STD_LOGIC;
                 signal ap_cpu_jtag_debug_module_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal ap_cpu_jtag_debug_module_resetrequest : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal ap_cpu_data_master_granted_ap_cpu_jtag_debug_module : OUT STD_LOGIC;
                 signal ap_cpu_data_master_qualified_request_ap_cpu_jtag_debug_module : OUT STD_LOGIC;
                 signal ap_cpu_data_master_read_data_valid_ap_cpu_jtag_debug_module : OUT STD_LOGIC;
                 signal ap_cpu_data_master_requests_ap_cpu_jtag_debug_module : OUT STD_LOGIC;
                 signal ap_cpu_instruction_master_granted_ap_cpu_jtag_debug_module : OUT STD_LOGIC;
                 signal ap_cpu_instruction_master_qualified_request_ap_cpu_jtag_debug_module : OUT STD_LOGIC;
                 signal ap_cpu_instruction_master_read_data_valid_ap_cpu_jtag_debug_module : OUT STD_LOGIC;
                 signal ap_cpu_instruction_master_requests_ap_cpu_jtag_debug_module : OUT STD_LOGIC;
                 signal ap_cpu_jtag_debug_module_address : OUT STD_LOGIC_VECTOR (8 DOWNTO 0);
                 signal ap_cpu_jtag_debug_module_begintransfer : OUT STD_LOGIC;
                 signal ap_cpu_jtag_debug_module_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal ap_cpu_jtag_debug_module_chipselect : OUT STD_LOGIC;
                 signal ap_cpu_jtag_debug_module_debugaccess : OUT STD_LOGIC;
                 signal ap_cpu_jtag_debug_module_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal ap_cpu_jtag_debug_module_reset_n : OUT STD_LOGIC;
                 signal ap_cpu_jtag_debug_module_resetrequest_from_sa : OUT STD_LOGIC;
                 signal ap_cpu_jtag_debug_module_write : OUT STD_LOGIC;
                 signal ap_cpu_jtag_debug_module_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal d1_ap_cpu_jtag_debug_module_end_xfer : OUT STD_LOGIC
              );
end entity ap_cpu_jtag_debug_module_arbitrator;


architecture europa of ap_cpu_jtag_debug_module_arbitrator is
                signal ap_cpu_data_master_arbiterlock :  STD_LOGIC;
                signal ap_cpu_data_master_arbiterlock2 :  STD_LOGIC;
                signal ap_cpu_data_master_continuerequest :  STD_LOGIC;
                signal ap_cpu_data_master_saved_grant_ap_cpu_jtag_debug_module :  STD_LOGIC;
                signal ap_cpu_instruction_master_arbiterlock :  STD_LOGIC;
                signal ap_cpu_instruction_master_arbiterlock2 :  STD_LOGIC;
                signal ap_cpu_instruction_master_continuerequest :  STD_LOGIC;
                signal ap_cpu_instruction_master_saved_grant_ap_cpu_jtag_debug_module :  STD_LOGIC;
                signal ap_cpu_jtag_debug_module_allgrants :  STD_LOGIC;
                signal ap_cpu_jtag_debug_module_allow_new_arb_cycle :  STD_LOGIC;
                signal ap_cpu_jtag_debug_module_any_bursting_master_saved_grant :  STD_LOGIC;
                signal ap_cpu_jtag_debug_module_any_continuerequest :  STD_LOGIC;
                signal ap_cpu_jtag_debug_module_arb_addend :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal ap_cpu_jtag_debug_module_arb_counter_enable :  STD_LOGIC;
                signal ap_cpu_jtag_debug_module_arb_share_counter :  STD_LOGIC;
                signal ap_cpu_jtag_debug_module_arb_share_counter_next_value :  STD_LOGIC;
                signal ap_cpu_jtag_debug_module_arb_share_set_values :  STD_LOGIC;
                signal ap_cpu_jtag_debug_module_arb_winner :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal ap_cpu_jtag_debug_module_arbitration_holdoff_internal :  STD_LOGIC;
                signal ap_cpu_jtag_debug_module_beginbursttransfer_internal :  STD_LOGIC;
                signal ap_cpu_jtag_debug_module_begins_xfer :  STD_LOGIC;
                signal ap_cpu_jtag_debug_module_chosen_master_double_vector :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal ap_cpu_jtag_debug_module_chosen_master_rot_left :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal ap_cpu_jtag_debug_module_end_xfer :  STD_LOGIC;
                signal ap_cpu_jtag_debug_module_firsttransfer :  STD_LOGIC;
                signal ap_cpu_jtag_debug_module_grant_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal ap_cpu_jtag_debug_module_in_a_read_cycle :  STD_LOGIC;
                signal ap_cpu_jtag_debug_module_in_a_write_cycle :  STD_LOGIC;
                signal ap_cpu_jtag_debug_module_master_qreq_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal ap_cpu_jtag_debug_module_non_bursting_master_requests :  STD_LOGIC;
                signal ap_cpu_jtag_debug_module_reg_firsttransfer :  STD_LOGIC;
                signal ap_cpu_jtag_debug_module_saved_chosen_master_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal ap_cpu_jtag_debug_module_slavearbiterlockenable :  STD_LOGIC;
                signal ap_cpu_jtag_debug_module_slavearbiterlockenable2 :  STD_LOGIC;
                signal ap_cpu_jtag_debug_module_unreg_firsttransfer :  STD_LOGIC;
                signal ap_cpu_jtag_debug_module_waits_for_read :  STD_LOGIC;
                signal ap_cpu_jtag_debug_module_waits_for_write :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_ap_cpu_jtag_debug_module :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_ap_cpu_data_master_granted_ap_cpu_jtag_debug_module :  STD_LOGIC;
                signal internal_ap_cpu_data_master_qualified_request_ap_cpu_jtag_debug_module :  STD_LOGIC;
                signal internal_ap_cpu_data_master_requests_ap_cpu_jtag_debug_module :  STD_LOGIC;
                signal internal_ap_cpu_instruction_master_granted_ap_cpu_jtag_debug_module :  STD_LOGIC;
                signal internal_ap_cpu_instruction_master_qualified_request_ap_cpu_jtag_debug_module :  STD_LOGIC;
                signal internal_ap_cpu_instruction_master_requests_ap_cpu_jtag_debug_module :  STD_LOGIC;
                signal last_cycle_ap_cpu_data_master_granted_slave_ap_cpu_jtag_debug_module :  STD_LOGIC;
                signal last_cycle_ap_cpu_instruction_master_granted_slave_ap_cpu_jtag_debug_module :  STD_LOGIC;
                signal shifted_address_to_ap_cpu_jtag_debug_module_from_ap_cpu_data_master :  STD_LOGIC_VECTOR (25 DOWNTO 0);
                signal shifted_address_to_ap_cpu_jtag_debug_module_from_ap_cpu_instruction_master :  STD_LOGIC_VECTOR (25 DOWNTO 0);
                signal wait_for_ap_cpu_jtag_debug_module_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT ap_cpu_jtag_debug_module_end_xfer;
    end if;

  end process;

  ap_cpu_jtag_debug_module_begins_xfer <= NOT d1_reasons_to_wait AND ((internal_ap_cpu_data_master_qualified_request_ap_cpu_jtag_debug_module OR internal_ap_cpu_instruction_master_qualified_request_ap_cpu_jtag_debug_module));
  --assign ap_cpu_jtag_debug_module_readdata_from_sa = ap_cpu_jtag_debug_module_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  ap_cpu_jtag_debug_module_readdata_from_sa <= ap_cpu_jtag_debug_module_readdata;
  internal_ap_cpu_data_master_requests_ap_cpu_jtag_debug_module <= to_std_logic(((Std_Logic_Vector'(ap_cpu_data_master_address_to_slave(25 DOWNTO 11) & std_logic_vector'("00000000000")) = std_logic_vector'("11000000100000100000000000")))) AND ((ap_cpu_data_master_read OR ap_cpu_data_master_write));
  --ap_cpu_jtag_debug_module_arb_share_counter set values, which is an e_mux
  ap_cpu_jtag_debug_module_arb_share_set_values <= std_logic'('1');
  --ap_cpu_jtag_debug_module_non_bursting_master_requests mux, which is an e_mux
  ap_cpu_jtag_debug_module_non_bursting_master_requests <= ((internal_ap_cpu_data_master_requests_ap_cpu_jtag_debug_module OR internal_ap_cpu_instruction_master_requests_ap_cpu_jtag_debug_module) OR internal_ap_cpu_data_master_requests_ap_cpu_jtag_debug_module) OR internal_ap_cpu_instruction_master_requests_ap_cpu_jtag_debug_module;
  --ap_cpu_jtag_debug_module_any_bursting_master_saved_grant mux, which is an e_mux
  ap_cpu_jtag_debug_module_any_bursting_master_saved_grant <= std_logic'('0');
  --ap_cpu_jtag_debug_module_arb_share_counter_next_value assignment, which is an e_assign
  ap_cpu_jtag_debug_module_arb_share_counter_next_value <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(ap_cpu_jtag_debug_module_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(ap_cpu_jtag_debug_module_arb_share_set_values))) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(ap_cpu_jtag_debug_module_arb_share_counter) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(ap_cpu_jtag_debug_module_arb_share_counter))) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))));
  --ap_cpu_jtag_debug_module_allgrants all slave grants, which is an e_mux
  ap_cpu_jtag_debug_module_allgrants <= (((or_reduce(ap_cpu_jtag_debug_module_grant_vector)) OR (or_reduce(ap_cpu_jtag_debug_module_grant_vector))) OR (or_reduce(ap_cpu_jtag_debug_module_grant_vector))) OR (or_reduce(ap_cpu_jtag_debug_module_grant_vector));
  --ap_cpu_jtag_debug_module_end_xfer assignment, which is an e_assign
  ap_cpu_jtag_debug_module_end_xfer <= NOT ((ap_cpu_jtag_debug_module_waits_for_read OR ap_cpu_jtag_debug_module_waits_for_write));
  --end_xfer_arb_share_counter_term_ap_cpu_jtag_debug_module arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_ap_cpu_jtag_debug_module <= ap_cpu_jtag_debug_module_end_xfer AND (((NOT ap_cpu_jtag_debug_module_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --ap_cpu_jtag_debug_module_arb_share_counter arbitration counter enable, which is an e_assign
  ap_cpu_jtag_debug_module_arb_counter_enable <= ((end_xfer_arb_share_counter_term_ap_cpu_jtag_debug_module AND ap_cpu_jtag_debug_module_allgrants)) OR ((end_xfer_arb_share_counter_term_ap_cpu_jtag_debug_module AND NOT ap_cpu_jtag_debug_module_non_bursting_master_requests));
  --ap_cpu_jtag_debug_module_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      ap_cpu_jtag_debug_module_arb_share_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(ap_cpu_jtag_debug_module_arb_counter_enable) = '1' then 
        ap_cpu_jtag_debug_module_arb_share_counter <= ap_cpu_jtag_debug_module_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --ap_cpu_jtag_debug_module_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      ap_cpu_jtag_debug_module_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((or_reduce(ap_cpu_jtag_debug_module_master_qreq_vector) AND end_xfer_arb_share_counter_term_ap_cpu_jtag_debug_module)) OR ((end_xfer_arb_share_counter_term_ap_cpu_jtag_debug_module AND NOT ap_cpu_jtag_debug_module_non_bursting_master_requests)))) = '1' then 
        ap_cpu_jtag_debug_module_slavearbiterlockenable <= ap_cpu_jtag_debug_module_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --ap_cpu/data_master ap_cpu/jtag_debug_module arbiterlock, which is an e_assign
  ap_cpu_data_master_arbiterlock <= ap_cpu_jtag_debug_module_slavearbiterlockenable AND ap_cpu_data_master_continuerequest;
  --ap_cpu_jtag_debug_module_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  ap_cpu_jtag_debug_module_slavearbiterlockenable2 <= ap_cpu_jtag_debug_module_arb_share_counter_next_value;
  --ap_cpu/data_master ap_cpu/jtag_debug_module arbiterlock2, which is an e_assign
  ap_cpu_data_master_arbiterlock2 <= ap_cpu_jtag_debug_module_slavearbiterlockenable2 AND ap_cpu_data_master_continuerequest;
  --ap_cpu/instruction_master ap_cpu/jtag_debug_module arbiterlock, which is an e_assign
  ap_cpu_instruction_master_arbiterlock <= ap_cpu_jtag_debug_module_slavearbiterlockenable AND ap_cpu_instruction_master_continuerequest;
  --ap_cpu/instruction_master ap_cpu/jtag_debug_module arbiterlock2, which is an e_assign
  ap_cpu_instruction_master_arbiterlock2 <= ap_cpu_jtag_debug_module_slavearbiterlockenable2 AND ap_cpu_instruction_master_continuerequest;
  --ap_cpu/instruction_master granted ap_cpu/jtag_debug_module last time, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      last_cycle_ap_cpu_instruction_master_granted_slave_ap_cpu_jtag_debug_module <= std_logic'('0');
    elsif clk'event and clk = '1' then
      last_cycle_ap_cpu_instruction_master_granted_slave_ap_cpu_jtag_debug_module <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(ap_cpu_instruction_master_saved_grant_ap_cpu_jtag_debug_module) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((ap_cpu_jtag_debug_module_arbitration_holdoff_internal OR NOT internal_ap_cpu_instruction_master_requests_ap_cpu_jtag_debug_module))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_ap_cpu_instruction_master_granted_slave_ap_cpu_jtag_debug_module))))));
    end if;

  end process;

  --ap_cpu_instruction_master_continuerequest continued request, which is an e_mux
  ap_cpu_instruction_master_continuerequest <= last_cycle_ap_cpu_instruction_master_granted_slave_ap_cpu_jtag_debug_module AND internal_ap_cpu_instruction_master_requests_ap_cpu_jtag_debug_module;
  --ap_cpu_jtag_debug_module_any_continuerequest at least one master continues requesting, which is an e_mux
  ap_cpu_jtag_debug_module_any_continuerequest <= ap_cpu_instruction_master_continuerequest OR ap_cpu_data_master_continuerequest;
  internal_ap_cpu_data_master_qualified_request_ap_cpu_jtag_debug_module <= internal_ap_cpu_data_master_requests_ap_cpu_jtag_debug_module AND NOT (((((NOT ap_cpu_data_master_waitrequest) AND ap_cpu_data_master_write)) OR ap_cpu_instruction_master_arbiterlock));
  --ap_cpu_jtag_debug_module_writedata mux, which is an e_mux
  ap_cpu_jtag_debug_module_writedata <= ap_cpu_data_master_writedata;
  internal_ap_cpu_instruction_master_requests_ap_cpu_jtag_debug_module <= ((to_std_logic(((Std_Logic_Vector'(ap_cpu_instruction_master_address_to_slave(25 DOWNTO 11) & std_logic_vector'("00000000000")) = std_logic_vector'("11000000100000100000000000")))) AND (ap_cpu_instruction_master_read))) AND ap_cpu_instruction_master_read;
  --ap_cpu/data_master granted ap_cpu/jtag_debug_module last time, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      last_cycle_ap_cpu_data_master_granted_slave_ap_cpu_jtag_debug_module <= std_logic'('0');
    elsif clk'event and clk = '1' then
      last_cycle_ap_cpu_data_master_granted_slave_ap_cpu_jtag_debug_module <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(ap_cpu_data_master_saved_grant_ap_cpu_jtag_debug_module) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((ap_cpu_jtag_debug_module_arbitration_holdoff_internal OR NOT internal_ap_cpu_data_master_requests_ap_cpu_jtag_debug_module))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_ap_cpu_data_master_granted_slave_ap_cpu_jtag_debug_module))))));
    end if;

  end process;

  --ap_cpu_data_master_continuerequest continued request, which is an e_mux
  ap_cpu_data_master_continuerequest <= last_cycle_ap_cpu_data_master_granted_slave_ap_cpu_jtag_debug_module AND internal_ap_cpu_data_master_requests_ap_cpu_jtag_debug_module;
  internal_ap_cpu_instruction_master_qualified_request_ap_cpu_jtag_debug_module <= internal_ap_cpu_instruction_master_requests_ap_cpu_jtag_debug_module AND NOT ((((ap_cpu_instruction_master_read AND ((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(ap_cpu_instruction_master_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000")))) OR (ap_cpu_instruction_master_read_data_valid_sdram_0_s1_shift_register))))) OR ap_cpu_data_master_arbiterlock));
  --local readdatavalid ap_cpu_instruction_master_read_data_valid_ap_cpu_jtag_debug_module, which is an e_mux
  ap_cpu_instruction_master_read_data_valid_ap_cpu_jtag_debug_module <= (internal_ap_cpu_instruction_master_granted_ap_cpu_jtag_debug_module AND ap_cpu_instruction_master_read) AND NOT ap_cpu_jtag_debug_module_waits_for_read;
  --allow new arb cycle for ap_cpu/jtag_debug_module, which is an e_assign
  ap_cpu_jtag_debug_module_allow_new_arb_cycle <= NOT ap_cpu_data_master_arbiterlock AND NOT ap_cpu_instruction_master_arbiterlock;
  --ap_cpu/instruction_master assignment into master qualified-requests vector for ap_cpu/jtag_debug_module, which is an e_assign
  ap_cpu_jtag_debug_module_master_qreq_vector(0) <= internal_ap_cpu_instruction_master_qualified_request_ap_cpu_jtag_debug_module;
  --ap_cpu/instruction_master grant ap_cpu/jtag_debug_module, which is an e_assign
  internal_ap_cpu_instruction_master_granted_ap_cpu_jtag_debug_module <= ap_cpu_jtag_debug_module_grant_vector(0);
  --ap_cpu/instruction_master saved-grant ap_cpu/jtag_debug_module, which is an e_assign
  ap_cpu_instruction_master_saved_grant_ap_cpu_jtag_debug_module <= ap_cpu_jtag_debug_module_arb_winner(0) AND internal_ap_cpu_instruction_master_requests_ap_cpu_jtag_debug_module;
  --ap_cpu/data_master assignment into master qualified-requests vector for ap_cpu/jtag_debug_module, which is an e_assign
  ap_cpu_jtag_debug_module_master_qreq_vector(1) <= internal_ap_cpu_data_master_qualified_request_ap_cpu_jtag_debug_module;
  --ap_cpu/data_master grant ap_cpu/jtag_debug_module, which is an e_assign
  internal_ap_cpu_data_master_granted_ap_cpu_jtag_debug_module <= ap_cpu_jtag_debug_module_grant_vector(1);
  --ap_cpu/data_master saved-grant ap_cpu/jtag_debug_module, which is an e_assign
  ap_cpu_data_master_saved_grant_ap_cpu_jtag_debug_module <= ap_cpu_jtag_debug_module_arb_winner(1) AND internal_ap_cpu_data_master_requests_ap_cpu_jtag_debug_module;
  --ap_cpu/jtag_debug_module chosen-master double-vector, which is an e_assign
  ap_cpu_jtag_debug_module_chosen_master_double_vector <= A_EXT (((std_logic_vector'("0") & ((ap_cpu_jtag_debug_module_master_qreq_vector & ap_cpu_jtag_debug_module_master_qreq_vector))) AND (((std_logic_vector'("0") & (Std_Logic_Vector'(NOT ap_cpu_jtag_debug_module_master_qreq_vector & NOT ap_cpu_jtag_debug_module_master_qreq_vector))) + (std_logic_vector'("000") & (ap_cpu_jtag_debug_module_arb_addend))))), 4);
  --stable onehot encoding of arb winner
  ap_cpu_jtag_debug_module_arb_winner <= A_WE_StdLogicVector((std_logic'(((ap_cpu_jtag_debug_module_allow_new_arb_cycle AND or_reduce(ap_cpu_jtag_debug_module_grant_vector)))) = '1'), ap_cpu_jtag_debug_module_grant_vector, ap_cpu_jtag_debug_module_saved_chosen_master_vector);
  --saved ap_cpu_jtag_debug_module_grant_vector, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      ap_cpu_jtag_debug_module_saved_chosen_master_vector <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      if std_logic'(ap_cpu_jtag_debug_module_allow_new_arb_cycle) = '1' then 
        ap_cpu_jtag_debug_module_saved_chosen_master_vector <= A_WE_StdLogicVector((std_logic'(or_reduce(ap_cpu_jtag_debug_module_grant_vector)) = '1'), ap_cpu_jtag_debug_module_grant_vector, ap_cpu_jtag_debug_module_saved_chosen_master_vector);
      end if;
    end if;

  end process;

  --onehot encoding of chosen master
  ap_cpu_jtag_debug_module_grant_vector <= Std_Logic_Vector'(A_ToStdLogicVector(((ap_cpu_jtag_debug_module_chosen_master_double_vector(1) OR ap_cpu_jtag_debug_module_chosen_master_double_vector(3)))) & A_ToStdLogicVector(((ap_cpu_jtag_debug_module_chosen_master_double_vector(0) OR ap_cpu_jtag_debug_module_chosen_master_double_vector(2)))));
  --ap_cpu/jtag_debug_module chosen master rotated left, which is an e_assign
  ap_cpu_jtag_debug_module_chosen_master_rot_left <= A_EXT (A_WE_StdLogicVector((((A_SLL(ap_cpu_jtag_debug_module_arb_winner,std_logic_vector'("00000000000000000000000000000001")))) /= std_logic_vector'("00")), (std_logic_vector'("000000000000000000000000000000") & ((A_SLL(ap_cpu_jtag_debug_module_arb_winner,std_logic_vector'("00000000000000000000000000000001"))))), std_logic_vector'("00000000000000000000000000000001")), 2);
  --ap_cpu/jtag_debug_module's addend for next-master-grant
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      ap_cpu_jtag_debug_module_arb_addend <= std_logic_vector'("01");
    elsif clk'event and clk = '1' then
      if std_logic'(or_reduce(ap_cpu_jtag_debug_module_grant_vector)) = '1' then 
        ap_cpu_jtag_debug_module_arb_addend <= A_WE_StdLogicVector((std_logic'(ap_cpu_jtag_debug_module_end_xfer) = '1'), ap_cpu_jtag_debug_module_chosen_master_rot_left, ap_cpu_jtag_debug_module_grant_vector);
      end if;
    end if;

  end process;

  ap_cpu_jtag_debug_module_begintransfer <= ap_cpu_jtag_debug_module_begins_xfer;
  --ap_cpu_jtag_debug_module_reset_n assignment, which is an e_assign
  ap_cpu_jtag_debug_module_reset_n <= reset_n;
  --assign ap_cpu_jtag_debug_module_resetrequest_from_sa = ap_cpu_jtag_debug_module_resetrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  ap_cpu_jtag_debug_module_resetrequest_from_sa <= ap_cpu_jtag_debug_module_resetrequest;
  ap_cpu_jtag_debug_module_chipselect <= internal_ap_cpu_data_master_granted_ap_cpu_jtag_debug_module OR internal_ap_cpu_instruction_master_granted_ap_cpu_jtag_debug_module;
  --ap_cpu_jtag_debug_module_firsttransfer first transaction, which is an e_assign
  ap_cpu_jtag_debug_module_firsttransfer <= A_WE_StdLogic((std_logic'(ap_cpu_jtag_debug_module_begins_xfer) = '1'), ap_cpu_jtag_debug_module_unreg_firsttransfer, ap_cpu_jtag_debug_module_reg_firsttransfer);
  --ap_cpu_jtag_debug_module_unreg_firsttransfer first transaction, which is an e_assign
  ap_cpu_jtag_debug_module_unreg_firsttransfer <= NOT ((ap_cpu_jtag_debug_module_slavearbiterlockenable AND ap_cpu_jtag_debug_module_any_continuerequest));
  --ap_cpu_jtag_debug_module_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      ap_cpu_jtag_debug_module_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(ap_cpu_jtag_debug_module_begins_xfer) = '1' then 
        ap_cpu_jtag_debug_module_reg_firsttransfer <= ap_cpu_jtag_debug_module_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --ap_cpu_jtag_debug_module_beginbursttransfer_internal begin burst transfer, which is an e_assign
  ap_cpu_jtag_debug_module_beginbursttransfer_internal <= ap_cpu_jtag_debug_module_begins_xfer;
  --ap_cpu_jtag_debug_module_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  ap_cpu_jtag_debug_module_arbitration_holdoff_internal <= ap_cpu_jtag_debug_module_begins_xfer AND ap_cpu_jtag_debug_module_firsttransfer;
  --ap_cpu_jtag_debug_module_write assignment, which is an e_mux
  ap_cpu_jtag_debug_module_write <= internal_ap_cpu_data_master_granted_ap_cpu_jtag_debug_module AND ap_cpu_data_master_write;
  shifted_address_to_ap_cpu_jtag_debug_module_from_ap_cpu_data_master <= ap_cpu_data_master_address_to_slave;
  --ap_cpu_jtag_debug_module_address mux, which is an e_mux
  ap_cpu_jtag_debug_module_address <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_ap_cpu_data_master_granted_ap_cpu_jtag_debug_module)) = '1'), (A_SRL(shifted_address_to_ap_cpu_jtag_debug_module_from_ap_cpu_data_master,std_logic_vector'("00000000000000000000000000000010"))), (A_SRL(shifted_address_to_ap_cpu_jtag_debug_module_from_ap_cpu_instruction_master,std_logic_vector'("00000000000000000000000000000010")))), 9);
  shifted_address_to_ap_cpu_jtag_debug_module_from_ap_cpu_instruction_master <= ap_cpu_instruction_master_address_to_slave;
  --d1_ap_cpu_jtag_debug_module_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_ap_cpu_jtag_debug_module_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_ap_cpu_jtag_debug_module_end_xfer <= ap_cpu_jtag_debug_module_end_xfer;
    end if;

  end process;

  --ap_cpu_jtag_debug_module_waits_for_read in a cycle, which is an e_mux
  ap_cpu_jtag_debug_module_waits_for_read <= ap_cpu_jtag_debug_module_in_a_read_cycle AND ap_cpu_jtag_debug_module_begins_xfer;
  --ap_cpu_jtag_debug_module_in_a_read_cycle assignment, which is an e_assign
  ap_cpu_jtag_debug_module_in_a_read_cycle <= ((internal_ap_cpu_data_master_granted_ap_cpu_jtag_debug_module AND ap_cpu_data_master_read)) OR ((internal_ap_cpu_instruction_master_granted_ap_cpu_jtag_debug_module AND ap_cpu_instruction_master_read));
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= ap_cpu_jtag_debug_module_in_a_read_cycle;
  --ap_cpu_jtag_debug_module_waits_for_write in a cycle, which is an e_mux
  ap_cpu_jtag_debug_module_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(ap_cpu_jtag_debug_module_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --ap_cpu_jtag_debug_module_in_a_write_cycle assignment, which is an e_assign
  ap_cpu_jtag_debug_module_in_a_write_cycle <= internal_ap_cpu_data_master_granted_ap_cpu_jtag_debug_module AND ap_cpu_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= ap_cpu_jtag_debug_module_in_a_write_cycle;
  wait_for_ap_cpu_jtag_debug_module_counter <= std_logic'('0');
  --ap_cpu_jtag_debug_module_byteenable byte enable port mux, which is an e_mux
  ap_cpu_jtag_debug_module_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_ap_cpu_data_master_granted_ap_cpu_jtag_debug_module)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (ap_cpu_data_master_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))), 4);
  --debugaccess mux, which is an e_mux
  ap_cpu_jtag_debug_module_debugaccess <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((internal_ap_cpu_data_master_granted_ap_cpu_jtag_debug_module)) = '1'), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(ap_cpu_data_master_debugaccess))), std_logic_vector'("00000000000000000000000000000000")));
  --vhdl renameroo for output signals
  ap_cpu_data_master_granted_ap_cpu_jtag_debug_module <= internal_ap_cpu_data_master_granted_ap_cpu_jtag_debug_module;
  --vhdl renameroo for output signals
  ap_cpu_data_master_qualified_request_ap_cpu_jtag_debug_module <= internal_ap_cpu_data_master_qualified_request_ap_cpu_jtag_debug_module;
  --vhdl renameroo for output signals
  ap_cpu_data_master_requests_ap_cpu_jtag_debug_module <= internal_ap_cpu_data_master_requests_ap_cpu_jtag_debug_module;
  --vhdl renameroo for output signals
  ap_cpu_instruction_master_granted_ap_cpu_jtag_debug_module <= internal_ap_cpu_instruction_master_granted_ap_cpu_jtag_debug_module;
  --vhdl renameroo for output signals
  ap_cpu_instruction_master_qualified_request_ap_cpu_jtag_debug_module <= internal_ap_cpu_instruction_master_qualified_request_ap_cpu_jtag_debug_module;
  --vhdl renameroo for output signals
  ap_cpu_instruction_master_requests_ap_cpu_jtag_debug_module <= internal_ap_cpu_instruction_master_requests_ap_cpu_jtag_debug_module;
--synthesis translate_off
    --ap_cpu/jtag_debug_module enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --grant signals are active simultaneously, which is an e_process
    process (clk)
    VARIABLE write_line : line;
    begin
      if clk'event and clk = '1' then
        if (std_logic_vector'("000000000000000000000000000000") & (((std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(internal_ap_cpu_data_master_granted_ap_cpu_jtag_debug_module))) + (std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(internal_ap_cpu_instruction_master_granted_ap_cpu_jtag_debug_module))))))>std_logic_vector'("00000000000000000000000000000001") then 
          write(write_line, now);
          write(write_line, string'(": "));
          write(write_line, string'("> 1 of grant signals are active simultaneously"));
          write(output, write_line.all);
          deallocate (write_line);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --saved_grant signals are active simultaneously, which is an e_process
    process (clk)
    VARIABLE write_line1 : line;
    begin
      if clk'event and clk = '1' then
        if (std_logic_vector'("000000000000000000000000000000") & (((std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(ap_cpu_data_master_saved_grant_ap_cpu_jtag_debug_module))) + (std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(ap_cpu_instruction_master_saved_grant_ap_cpu_jtag_debug_module))))))>std_logic_vector'("00000000000000000000000000000001") then 
          write(write_line1, now);
          write(write_line1, string'(": "));
          write(write_line1, string'("> 1 of saved_grant signals are active simultaneously"));
          write(output, write_line1.all);
          deallocate (write_line1);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity sync_irq_s1_irq_from_sa_clock_crossing_ap_cpu_data_master_module is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC
              );
end entity sync_irq_s1_irq_from_sa_clock_crossing_ap_cpu_data_master_module;


architecture europa of sync_irq_s1_irq_from_sa_clock_crossing_ap_cpu_data_master_module is
                signal data_in_d1 :  STD_LOGIC;
attribute ALTERA_ATTRIBUTE : string;
attribute ALTERA_ATTRIBUTE of data_in_d1 : signal is "{-from ""*""} CUT=ON ; PRESERVE_REGISTER=ON";
attribute ALTERA_ATTRIBUTE of data_out : signal is "PRESERVE_REGISTER=ON";

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      data_in_d1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      data_in_d1 <= data_in;
    end if;

  end process;

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      data_out <= std_logic'('0');
    elsif clk'event and clk = '1' then
      data_out <= data_in_d1;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity system_timer_ap_s1_irq_from_sa_clock_crossing_ap_cpu_data_master_module is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC
              );
end entity system_timer_ap_s1_irq_from_sa_clock_crossing_ap_cpu_data_master_module;


architecture europa of system_timer_ap_s1_irq_from_sa_clock_crossing_ap_cpu_data_master_module is
                signal data_in_d1 :  STD_LOGIC;
attribute ALTERA_ATTRIBUTE : string;
attribute ALTERA_ATTRIBUTE of data_in_d1 : signal is "{-from ""*""} CUT=ON ; PRESERVE_REGISTER=ON";
attribute ALTERA_ATTRIBUTE of data_out : signal is "PRESERVE_REGISTER=ON";

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      data_in_d1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      data_in_d1 <= data_in;
    end if;

  end process;

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      data_out <= std_logic'('0');
    elsif clk'event and clk = '1' then
      data_out <= data_in_d1;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity ap_cpu_data_master_arbitrator is 
        port (
              -- inputs:
                 signal ap_cpu_data_master_address : IN STD_LOGIC_VECTOR (25 DOWNTO 0);
                 signal ap_cpu_data_master_granted_ap_cpu_jtag_debug_module : IN STD_LOGIC;
                 signal ap_cpu_data_master_granted_clock_crossing_1_s1 : IN STD_LOGIC;
                 signal ap_cpu_data_master_granted_cnApi_Av2Av_0_ap : IN STD_LOGIC;
                 signal ap_cpu_data_master_granted_jtag_uart_1_avalon_jtag_slave : IN STD_LOGIC;
                 signal ap_cpu_data_master_granted_sdram_0_s1 : IN STD_LOGIC;
                 signal ap_cpu_data_master_qualified_request_ap_cpu_jtag_debug_module : IN STD_LOGIC;
                 signal ap_cpu_data_master_qualified_request_clock_crossing_1_s1 : IN STD_LOGIC;
                 signal ap_cpu_data_master_qualified_request_cnApi_Av2Av_0_ap : IN STD_LOGIC;
                 signal ap_cpu_data_master_qualified_request_jtag_uart_1_avalon_jtag_slave : IN STD_LOGIC;
                 signal ap_cpu_data_master_qualified_request_sdram_0_s1 : IN STD_LOGIC;
                 signal ap_cpu_data_master_read : IN STD_LOGIC;
                 signal ap_cpu_data_master_read_data_valid_ap_cpu_jtag_debug_module : IN STD_LOGIC;
                 signal ap_cpu_data_master_read_data_valid_clock_crossing_1_s1 : IN STD_LOGIC;
                 signal ap_cpu_data_master_read_data_valid_clock_crossing_1_s1_shift_register : IN STD_LOGIC;
                 signal ap_cpu_data_master_read_data_valid_cnApi_Av2Av_0_ap : IN STD_LOGIC;
                 signal ap_cpu_data_master_read_data_valid_jtag_uart_1_avalon_jtag_slave : IN STD_LOGIC;
                 signal ap_cpu_data_master_read_data_valid_sdram_0_s1 : IN STD_LOGIC;
                 signal ap_cpu_data_master_read_data_valid_sdram_0_s1_shift_register : IN STD_LOGIC;
                 signal ap_cpu_data_master_requests_ap_cpu_jtag_debug_module : IN STD_LOGIC;
                 signal ap_cpu_data_master_requests_clock_crossing_1_s1 : IN STD_LOGIC;
                 signal ap_cpu_data_master_requests_cnApi_Av2Av_0_ap : IN STD_LOGIC;
                 signal ap_cpu_data_master_requests_jtag_uart_1_avalon_jtag_slave : IN STD_LOGIC;
                 signal ap_cpu_data_master_requests_sdram_0_s1 : IN STD_LOGIC;
                 signal ap_cpu_data_master_write : IN STD_LOGIC;
                 signal ap_cpu_jtag_debug_module_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal clk : IN STD_LOGIC;
                 signal clk90Meg : IN STD_LOGIC;
                 signal clk90Meg_reset_n : IN STD_LOGIC;
                 signal clock_crossing_1_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal clock_crossing_1_s1_waitrequest_from_sa : IN STD_LOGIC;
                 signal cnApi_Av2Av_0_ap_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal cnApi_Av2Av_0_ap_wait_counter_eq_0 : IN STD_LOGIC;
                 signal d1_ap_cpu_jtag_debug_module_end_xfer : IN STD_LOGIC;
                 signal d1_clock_crossing_1_s1_end_xfer : IN STD_LOGIC;
                 signal d1_cnApi_Av2Av_0_ap_end_xfer : IN STD_LOGIC;
                 signal d1_jtag_uart_1_avalon_jtag_slave_end_xfer : IN STD_LOGIC;
                 signal d1_sdram_0_s1_end_xfer : IN STD_LOGIC;
                 signal jtag_uart_1_avalon_jtag_slave_irq_from_sa : IN STD_LOGIC;
                 signal jtag_uart_1_avalon_jtag_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal jtag_uart_1_avalon_jtag_slave_waitrequest_from_sa : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sdram_0_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal sdram_0_s1_waitrequest_from_sa : IN STD_LOGIC;
                 signal sync_irq_s1_irq_from_sa : IN STD_LOGIC;
                 signal system_timer_ap_s1_irq_from_sa : IN STD_LOGIC;

              -- outputs:
                 signal ap_cpu_data_master_address_to_slave : OUT STD_LOGIC_VECTOR (25 DOWNTO 0);
                 signal ap_cpu_data_master_irq : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal ap_cpu_data_master_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal ap_cpu_data_master_waitrequest : OUT STD_LOGIC
              );
end entity ap_cpu_data_master_arbitrator;


architecture europa of ap_cpu_data_master_arbitrator is
component sync_irq_s1_irq_from_sa_clock_crossing_ap_cpu_data_master_module is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC
                 );
end component sync_irq_s1_irq_from_sa_clock_crossing_ap_cpu_data_master_module;

component system_timer_ap_s1_irq_from_sa_clock_crossing_ap_cpu_data_master_module is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC
                 );
end component system_timer_ap_s1_irq_from_sa_clock_crossing_ap_cpu_data_master_module;

                signal ap_cpu_data_master_run :  STD_LOGIC;
                signal clk90Meg_sync_irq_s1_irq_from_sa :  STD_LOGIC;
                signal clk90Meg_system_timer_ap_s1_irq_from_sa :  STD_LOGIC;
                signal internal_ap_cpu_data_master_address_to_slave :  STD_LOGIC_VECTOR (25 DOWNTO 0);
                signal internal_ap_cpu_data_master_waitrequest :  STD_LOGIC;
                signal p1_registered_ap_cpu_data_master_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal r_0 :  STD_LOGIC;
                signal r_2 :  STD_LOGIC;
                signal registered_ap_cpu_data_master_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);

begin

  --r_0 master_run cascaded wait assignment, which is an e_assign
  r_0 <= Vector_To_Std_Logic(((((((((((((((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((ap_cpu_data_master_qualified_request_ap_cpu_jtag_debug_module OR NOT ap_cpu_data_master_requests_ap_cpu_jtag_debug_module)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((ap_cpu_data_master_granted_ap_cpu_jtag_debug_module OR NOT ap_cpu_data_master_qualified_request_ap_cpu_jtag_debug_module)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT ap_cpu_data_master_qualified_request_ap_cpu_jtag_debug_module OR NOT ap_cpu_data_master_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(ap_cpu_data_master_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT ap_cpu_data_master_qualified_request_ap_cpu_jtag_debug_module OR NOT ap_cpu_data_master_write)))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(ap_cpu_data_master_write)))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((ap_cpu_data_master_qualified_request_clock_crossing_1_s1 OR ap_cpu_data_master_read_data_valid_clock_crossing_1_s1) OR NOT ap_cpu_data_master_requests_clock_crossing_1_s1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((NOT ap_cpu_data_master_qualified_request_clock_crossing_1_s1 OR NOT ap_cpu_data_master_read) OR ((ap_cpu_data_master_read_data_valid_clock_crossing_1_s1 AND ap_cpu_data_master_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT ap_cpu_data_master_qualified_request_clock_crossing_1_s1 OR NOT ((ap_cpu_data_master_read OR ap_cpu_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT clock_crossing_1_s1_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((ap_cpu_data_master_read OR ap_cpu_data_master_write)))))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((ap_cpu_data_master_qualified_request_cnApi_Av2Av_0_ap OR NOT ap_cpu_data_master_requests_cnApi_Av2Av_0_ap)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT ap_cpu_data_master_qualified_request_cnApi_Av2Av_0_ap OR NOT ap_cpu_data_master_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT d1_cnApi_Av2Av_0_ap_end_xfer)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(ap_cpu_data_master_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT ap_cpu_data_master_qualified_request_cnApi_Av2Av_0_ap OR NOT ap_cpu_data_master_write)))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(ap_cpu_data_master_write)))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((ap_cpu_data_master_qualified_request_jtag_uart_1_avalon_jtag_slave OR NOT ap_cpu_data_master_requests_jtag_uart_1_avalon_jtag_slave)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT ap_cpu_data_master_qualified_request_jtag_uart_1_avalon_jtag_slave OR NOT ((ap_cpu_data_master_read OR ap_cpu_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT jtag_uart_1_avalon_jtag_slave_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((ap_cpu_data_master_read OR ap_cpu_data_master_write)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT ap_cpu_data_master_qualified_request_jtag_uart_1_avalon_jtag_slave OR NOT ((ap_cpu_data_master_read OR ap_cpu_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT jtag_uart_1_avalon_jtag_slave_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((ap_cpu_data_master_read OR ap_cpu_data_master_write)))))))))));
  --cascaded wait assignment, which is an e_assign
  ap_cpu_data_master_run <= r_0 AND r_2;
  --r_2 master_run cascaded wait assignment, which is an e_assign
  r_2 <= Vector_To_Std_Logic(((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((ap_cpu_data_master_qualified_request_sdram_0_s1 OR ap_cpu_data_master_read_data_valid_sdram_0_s1) OR NOT ap_cpu_data_master_requests_sdram_0_s1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((ap_cpu_data_master_granted_sdram_0_s1 OR NOT ap_cpu_data_master_qualified_request_sdram_0_s1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((NOT ap_cpu_data_master_qualified_request_sdram_0_s1 OR NOT ap_cpu_data_master_read) OR ((ap_cpu_data_master_read_data_valid_sdram_0_s1 AND ap_cpu_data_master_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT ap_cpu_data_master_qualified_request_sdram_0_s1 OR NOT ((ap_cpu_data_master_read OR ap_cpu_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT sdram_0_s1_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((ap_cpu_data_master_read OR ap_cpu_data_master_write)))))))))));
  --optimize select-logic by passing only those address bits which matter.
  internal_ap_cpu_data_master_address_to_slave <= ap_cpu_data_master_address(25 DOWNTO 0);
  --ap_cpu/data_master readdata mux, which is an e_mux
  ap_cpu_data_master_readdata <= (((((A_REP(NOT ap_cpu_data_master_requests_ap_cpu_jtag_debug_module, 32) OR ap_cpu_jtag_debug_module_readdata_from_sa)) AND ((A_REP(NOT ap_cpu_data_master_requests_clock_crossing_1_s1, 32) OR registered_ap_cpu_data_master_readdata))) AND ((A_REP(NOT ap_cpu_data_master_requests_cnApi_Av2Av_0_ap, 32) OR cnApi_Av2Av_0_ap_readdata_from_sa))) AND ((A_REP(NOT ap_cpu_data_master_requests_jtag_uart_1_avalon_jtag_slave, 32) OR registered_ap_cpu_data_master_readdata))) AND ((A_REP(NOT ap_cpu_data_master_requests_sdram_0_s1, 32) OR registered_ap_cpu_data_master_readdata));
  --actual waitrequest port, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      internal_ap_cpu_data_master_waitrequest <= Vector_To_Std_Logic(NOT std_logic_vector'("00000000000000000000000000000000"));
    elsif clk'event and clk = '1' then
      internal_ap_cpu_data_master_waitrequest <= Vector_To_Std_Logic(NOT (A_WE_StdLogicVector((std_logic'((NOT ((ap_cpu_data_master_read OR ap_cpu_data_master_write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((ap_cpu_data_master_run AND internal_ap_cpu_data_master_waitrequest))))))));
    end if;

  end process;

  --unpredictable registered wait state incoming data, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      registered_ap_cpu_data_master_readdata <= std_logic_vector'("00000000000000000000000000000000");
    elsif clk'event and clk = '1' then
      registered_ap_cpu_data_master_readdata <= p1_registered_ap_cpu_data_master_readdata;
    end if;

  end process;

  --registered readdata mux, which is an e_mux
  p1_registered_ap_cpu_data_master_readdata <= (((A_REP(NOT ap_cpu_data_master_requests_clock_crossing_1_s1, 32) OR clock_crossing_1_s1_readdata_from_sa)) AND ((A_REP(NOT ap_cpu_data_master_requests_jtag_uart_1_avalon_jtag_slave, 32) OR jtag_uart_1_avalon_jtag_slave_readdata_from_sa))) AND ((A_REP(NOT ap_cpu_data_master_requests_sdram_0_s1, 32) OR sdram_0_s1_readdata_from_sa));
  --irq assign, which is an e_assign
  ap_cpu_data_master_irq <= Std_Logic_Vector'(A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(jtag_uart_1_avalon_jtag_slave_irq_from_sa) & A_ToStdLogicVector(clk90Meg_system_timer_ap_s1_irq_from_sa) & A_ToStdLogicVector(clk90Meg_sync_irq_s1_irq_from_sa) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')));
  --sync_irq_s1_irq_from_sa from clk50Meg to clk90Meg
  sync_irq_s1_irq_from_sa_clock_crossing_ap_cpu_data_master : sync_irq_s1_irq_from_sa_clock_crossing_ap_cpu_data_master_module
    port map(
      data_out => clk90Meg_sync_irq_s1_irq_from_sa,
      clk => clk90Meg,
      data_in => sync_irq_s1_irq_from_sa,
      reset_n => clk90Meg_reset_n
    );


  --system_timer_ap_s1_irq_from_sa from clk50Meg to clk90Meg
  system_timer_ap_s1_irq_from_sa_clock_crossing_ap_cpu_data_master : system_timer_ap_s1_irq_from_sa_clock_crossing_ap_cpu_data_master_module
    port map(
      data_out => clk90Meg_system_timer_ap_s1_irq_from_sa,
      clk => clk90Meg,
      data_in => system_timer_ap_s1_irq_from_sa,
      reset_n => clk90Meg_reset_n
    );


  --vhdl renameroo for output signals
  ap_cpu_data_master_address_to_slave <= internal_ap_cpu_data_master_address_to_slave;
  --vhdl renameroo for output signals
  ap_cpu_data_master_waitrequest <= internal_ap_cpu_data_master_waitrequest;

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity ap_cpu_instruction_master_arbitrator is 
        port (
              -- inputs:
                 signal ap_cpu_instruction_master_address : IN STD_LOGIC_VECTOR (25 DOWNTO 0);
                 signal ap_cpu_instruction_master_granted_ap_cpu_jtag_debug_module : IN STD_LOGIC;
                 signal ap_cpu_instruction_master_granted_sdram_0_s1 : IN STD_LOGIC;
                 signal ap_cpu_instruction_master_qualified_request_ap_cpu_jtag_debug_module : IN STD_LOGIC;
                 signal ap_cpu_instruction_master_qualified_request_sdram_0_s1 : IN STD_LOGIC;
                 signal ap_cpu_instruction_master_read : IN STD_LOGIC;
                 signal ap_cpu_instruction_master_read_data_valid_ap_cpu_jtag_debug_module : IN STD_LOGIC;
                 signal ap_cpu_instruction_master_read_data_valid_sdram_0_s1 : IN STD_LOGIC;
                 signal ap_cpu_instruction_master_read_data_valid_sdram_0_s1_shift_register : IN STD_LOGIC;
                 signal ap_cpu_instruction_master_requests_ap_cpu_jtag_debug_module : IN STD_LOGIC;
                 signal ap_cpu_instruction_master_requests_sdram_0_s1 : IN STD_LOGIC;
                 signal ap_cpu_jtag_debug_module_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal clk : IN STD_LOGIC;
                 signal d1_ap_cpu_jtag_debug_module_end_xfer : IN STD_LOGIC;
                 signal d1_sdram_0_s1_end_xfer : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sdram_0_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal sdram_0_s1_waitrequest_from_sa : IN STD_LOGIC;

              -- outputs:
                 signal ap_cpu_instruction_master_address_to_slave : OUT STD_LOGIC_VECTOR (25 DOWNTO 0);
                 signal ap_cpu_instruction_master_latency_counter : OUT STD_LOGIC;
                 signal ap_cpu_instruction_master_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal ap_cpu_instruction_master_readdatavalid : OUT STD_LOGIC;
                 signal ap_cpu_instruction_master_waitrequest : OUT STD_LOGIC
              );
end entity ap_cpu_instruction_master_arbitrator;


architecture europa of ap_cpu_instruction_master_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal ap_cpu_instruction_master_address_last_time :  STD_LOGIC_VECTOR (25 DOWNTO 0);
                signal ap_cpu_instruction_master_is_granted_some_slave :  STD_LOGIC;
                signal ap_cpu_instruction_master_read_but_no_slave_selected :  STD_LOGIC;
                signal ap_cpu_instruction_master_read_last_time :  STD_LOGIC;
                signal ap_cpu_instruction_master_run :  STD_LOGIC;
                signal internal_ap_cpu_instruction_master_address_to_slave :  STD_LOGIC_VECTOR (25 DOWNTO 0);
                signal internal_ap_cpu_instruction_master_latency_counter :  STD_LOGIC;
                signal internal_ap_cpu_instruction_master_waitrequest :  STD_LOGIC;
                signal latency_load_value :  STD_LOGIC;
                signal p1_ap_cpu_instruction_master_latency_counter :  STD_LOGIC;
                signal pre_flush_ap_cpu_instruction_master_readdatavalid :  STD_LOGIC;
                signal r_0 :  STD_LOGIC;
                signal r_2 :  STD_LOGIC;

begin

  --r_0 master_run cascaded wait assignment, which is an e_assign
  r_0 <= Vector_To_Std_Logic((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((ap_cpu_instruction_master_qualified_request_ap_cpu_jtag_debug_module OR NOT ap_cpu_instruction_master_requests_ap_cpu_jtag_debug_module)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((ap_cpu_instruction_master_granted_ap_cpu_jtag_debug_module OR NOT ap_cpu_instruction_master_qualified_request_ap_cpu_jtag_debug_module)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT ap_cpu_instruction_master_qualified_request_ap_cpu_jtag_debug_module OR NOT ap_cpu_instruction_master_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT d1_ap_cpu_jtag_debug_module_end_xfer)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(ap_cpu_instruction_master_read)))))))));
  --cascaded wait assignment, which is an e_assign
  ap_cpu_instruction_master_run <= r_0 AND r_2;
  --r_2 master_run cascaded wait assignment, which is an e_assign
  r_2 <= Vector_To_Std_Logic((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((ap_cpu_instruction_master_qualified_request_sdram_0_s1 OR NOT ap_cpu_instruction_master_requests_sdram_0_s1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((ap_cpu_instruction_master_granted_sdram_0_s1 OR NOT ap_cpu_instruction_master_qualified_request_sdram_0_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT ap_cpu_instruction_master_qualified_request_sdram_0_s1 OR NOT ap_cpu_instruction_master_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT sdram_0_s1_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(ap_cpu_instruction_master_read)))))))));
  --optimize select-logic by passing only those address bits which matter.
  internal_ap_cpu_instruction_master_address_to_slave <= Std_Logic_Vector'(A_ToStdLogicVector(std_logic'('1')) & ap_cpu_instruction_master_address(24 DOWNTO 0));
  --ap_cpu_instruction_master_read_but_no_slave_selected assignment, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      ap_cpu_instruction_master_read_but_no_slave_selected <= std_logic'('0');
    elsif clk'event and clk = '1' then
      ap_cpu_instruction_master_read_but_no_slave_selected <= (ap_cpu_instruction_master_read AND ap_cpu_instruction_master_run) AND NOT ap_cpu_instruction_master_is_granted_some_slave;
    end if;

  end process;

  --some slave is getting selected, which is an e_mux
  ap_cpu_instruction_master_is_granted_some_slave <= ap_cpu_instruction_master_granted_ap_cpu_jtag_debug_module OR ap_cpu_instruction_master_granted_sdram_0_s1;
  --latent slave read data valids which may be flushed, which is an e_mux
  pre_flush_ap_cpu_instruction_master_readdatavalid <= ap_cpu_instruction_master_read_data_valid_sdram_0_s1;
  --latent slave read data valid which is not flushed, which is an e_mux
  ap_cpu_instruction_master_readdatavalid <= (((ap_cpu_instruction_master_read_but_no_slave_selected OR pre_flush_ap_cpu_instruction_master_readdatavalid) OR ap_cpu_instruction_master_read_data_valid_ap_cpu_jtag_debug_module) OR ap_cpu_instruction_master_read_but_no_slave_selected) OR pre_flush_ap_cpu_instruction_master_readdatavalid;
  --ap_cpu/instruction_master readdata mux, which is an e_mux
  ap_cpu_instruction_master_readdata <= ((A_REP(NOT ((ap_cpu_instruction_master_qualified_request_ap_cpu_jtag_debug_module AND ap_cpu_instruction_master_read)) , 32) OR ap_cpu_jtag_debug_module_readdata_from_sa)) AND ((A_REP(NOT ap_cpu_instruction_master_read_data_valid_sdram_0_s1, 32) OR sdram_0_s1_readdata_from_sa));
  --actual waitrequest port, which is an e_assign
  internal_ap_cpu_instruction_master_waitrequest <= NOT ap_cpu_instruction_master_run;
  --latent max counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      internal_ap_cpu_instruction_master_latency_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      internal_ap_cpu_instruction_master_latency_counter <= p1_ap_cpu_instruction_master_latency_counter;
    end if;

  end process;

  --latency counter load mux, which is an e_mux
  p1_ap_cpu_instruction_master_latency_counter <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(((ap_cpu_instruction_master_run AND ap_cpu_instruction_master_read))) = '1'), (std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(latency_load_value))), A_WE_StdLogicVector((std_logic'((internal_ap_cpu_instruction_master_latency_counter)) = '1'), ((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(internal_ap_cpu_instruction_master_latency_counter))) - std_logic_vector'("000000000000000000000000000000001")), std_logic_vector'("000000000000000000000000000000000"))));
  --read latency load values, which is an e_mux
  latency_load_value <= std_logic'('0');
  --vhdl renameroo for output signals
  ap_cpu_instruction_master_address_to_slave <= internal_ap_cpu_instruction_master_address_to_slave;
  --vhdl renameroo for output signals
  ap_cpu_instruction_master_latency_counter <= internal_ap_cpu_instruction_master_latency_counter;
  --vhdl renameroo for output signals
  ap_cpu_instruction_master_waitrequest <= internal_ap_cpu_instruction_master_waitrequest;
--synthesis translate_off
    --ap_cpu_instruction_master_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        ap_cpu_instruction_master_address_last_time <= std_logic_vector'("00000000000000000000000000");
      elsif clk'event and clk = '1' then
        ap_cpu_instruction_master_address_last_time <= ap_cpu_instruction_master_address;
      end if;

    end process;

    --ap_cpu/instruction_master waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_ap_cpu_instruction_master_waitrequest AND (ap_cpu_instruction_master_read);
      end if;

    end process;

    --ap_cpu_instruction_master_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line2 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((ap_cpu_instruction_master_address /= ap_cpu_instruction_master_address_last_time))))) = '1' then 
          write(write_line2, now);
          write(write_line2, string'(": "));
          write(write_line2, string'("ap_cpu_instruction_master_address did not heed wait!!!"));
          write(output, write_line2.all);
          deallocate (write_line2);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --ap_cpu_instruction_master_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        ap_cpu_instruction_master_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        ap_cpu_instruction_master_read_last_time <= ap_cpu_instruction_master_read;
      end if;

    end process;

    --ap_cpu_instruction_master_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line3 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(ap_cpu_instruction_master_read) /= std_logic'(ap_cpu_instruction_master_read_last_time)))))) = '1' then 
          write(write_line3, now);
          write(write_line3, string'(": "));
          write(write_line3, string'("ap_cpu_instruction_master_read did not heed wait!!!"));
          write(output, write_line3.all);
          deallocate (write_line3);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity button_pio_s1_arbitrator is 
        port (
              -- inputs:
                 signal button_pio_s1_readdata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal clk : IN STD_LOGIC;
                 signal clock_crossing_0_m1_address_to_slave : IN STD_LOGIC_VECTOR (6 DOWNTO 0);
                 signal clock_crossing_0_m1_latency_counter : IN STD_LOGIC;
                 signal clock_crossing_0_m1_nativeaddress : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
                 signal clock_crossing_0_m1_read : IN STD_LOGIC;
                 signal clock_crossing_0_m1_write : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal button_pio_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal button_pio_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal button_pio_s1_reset_n : OUT STD_LOGIC;
                 signal clock_crossing_0_m1_granted_button_pio_s1 : OUT STD_LOGIC;
                 signal clock_crossing_0_m1_qualified_request_button_pio_s1 : OUT STD_LOGIC;
                 signal clock_crossing_0_m1_read_data_valid_button_pio_s1 : OUT STD_LOGIC;
                 signal clock_crossing_0_m1_requests_button_pio_s1 : OUT STD_LOGIC;
                 signal d1_button_pio_s1_end_xfer : OUT STD_LOGIC
              );
end entity button_pio_s1_arbitrator;


architecture europa of button_pio_s1_arbitrator is
                signal button_pio_s1_allgrants :  STD_LOGIC;
                signal button_pio_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal button_pio_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal button_pio_s1_any_continuerequest :  STD_LOGIC;
                signal button_pio_s1_arb_counter_enable :  STD_LOGIC;
                signal button_pio_s1_arb_share_counter :  STD_LOGIC;
                signal button_pio_s1_arb_share_counter_next_value :  STD_LOGIC;
                signal button_pio_s1_arb_share_set_values :  STD_LOGIC;
                signal button_pio_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal button_pio_s1_begins_xfer :  STD_LOGIC;
                signal button_pio_s1_end_xfer :  STD_LOGIC;
                signal button_pio_s1_firsttransfer :  STD_LOGIC;
                signal button_pio_s1_grant_vector :  STD_LOGIC;
                signal button_pio_s1_in_a_read_cycle :  STD_LOGIC;
                signal button_pio_s1_in_a_write_cycle :  STD_LOGIC;
                signal button_pio_s1_master_qreq_vector :  STD_LOGIC;
                signal button_pio_s1_non_bursting_master_requests :  STD_LOGIC;
                signal button_pio_s1_reg_firsttransfer :  STD_LOGIC;
                signal button_pio_s1_slavearbiterlockenable :  STD_LOGIC;
                signal button_pio_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal button_pio_s1_unreg_firsttransfer :  STD_LOGIC;
                signal button_pio_s1_waits_for_read :  STD_LOGIC;
                signal button_pio_s1_waits_for_write :  STD_LOGIC;
                signal clock_crossing_0_m1_arbiterlock :  STD_LOGIC;
                signal clock_crossing_0_m1_arbiterlock2 :  STD_LOGIC;
                signal clock_crossing_0_m1_continuerequest :  STD_LOGIC;
                signal clock_crossing_0_m1_saved_grant_button_pio_s1 :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_button_pio_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_clock_crossing_0_m1_granted_button_pio_s1 :  STD_LOGIC;
                signal internal_clock_crossing_0_m1_qualified_request_button_pio_s1 :  STD_LOGIC;
                signal internal_clock_crossing_0_m1_requests_button_pio_s1 :  STD_LOGIC;
                signal wait_for_button_pio_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT button_pio_s1_end_xfer;
    end if;

  end process;

  button_pio_s1_begins_xfer <= NOT d1_reasons_to_wait AND (internal_clock_crossing_0_m1_qualified_request_button_pio_s1);
  --assign button_pio_s1_readdata_from_sa = button_pio_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  button_pio_s1_readdata_from_sa <= button_pio_s1_readdata;
  internal_clock_crossing_0_m1_requests_button_pio_s1 <= ((to_std_logic(((Std_Logic_Vector'(clock_crossing_0_m1_address_to_slave(6 DOWNTO 4) & std_logic_vector'("0000")) = std_logic_vector'("1010000")))) AND ((clock_crossing_0_m1_read OR clock_crossing_0_m1_write)))) AND clock_crossing_0_m1_read;
  --button_pio_s1_arb_share_counter set values, which is an e_mux
  button_pio_s1_arb_share_set_values <= std_logic'('1');
  --button_pio_s1_non_bursting_master_requests mux, which is an e_mux
  button_pio_s1_non_bursting_master_requests <= internal_clock_crossing_0_m1_requests_button_pio_s1;
  --button_pio_s1_any_bursting_master_saved_grant mux, which is an e_mux
  button_pio_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --button_pio_s1_arb_share_counter_next_value assignment, which is an e_assign
  button_pio_s1_arb_share_counter_next_value <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(button_pio_s1_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(button_pio_s1_arb_share_set_values))) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(button_pio_s1_arb_share_counter) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(button_pio_s1_arb_share_counter))) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))));
  --button_pio_s1_allgrants all slave grants, which is an e_mux
  button_pio_s1_allgrants <= button_pio_s1_grant_vector;
  --button_pio_s1_end_xfer assignment, which is an e_assign
  button_pio_s1_end_xfer <= NOT ((button_pio_s1_waits_for_read OR button_pio_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_button_pio_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_button_pio_s1 <= button_pio_s1_end_xfer AND (((NOT button_pio_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --button_pio_s1_arb_share_counter arbitration counter enable, which is an e_assign
  button_pio_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_button_pio_s1 AND button_pio_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_button_pio_s1 AND NOT button_pio_s1_non_bursting_master_requests));
  --button_pio_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      button_pio_s1_arb_share_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(button_pio_s1_arb_counter_enable) = '1' then 
        button_pio_s1_arb_share_counter <= button_pio_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --button_pio_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      button_pio_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((button_pio_s1_master_qreq_vector AND end_xfer_arb_share_counter_term_button_pio_s1)) OR ((end_xfer_arb_share_counter_term_button_pio_s1 AND NOT button_pio_s1_non_bursting_master_requests)))) = '1' then 
        button_pio_s1_slavearbiterlockenable <= button_pio_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --clock_crossing_0/m1 button_pio/s1 arbiterlock, which is an e_assign
  clock_crossing_0_m1_arbiterlock <= button_pio_s1_slavearbiterlockenable AND clock_crossing_0_m1_continuerequest;
  --button_pio_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  button_pio_s1_slavearbiterlockenable2 <= button_pio_s1_arb_share_counter_next_value;
  --clock_crossing_0/m1 button_pio/s1 arbiterlock2, which is an e_assign
  clock_crossing_0_m1_arbiterlock2 <= button_pio_s1_slavearbiterlockenable2 AND clock_crossing_0_m1_continuerequest;
  --button_pio_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  button_pio_s1_any_continuerequest <= std_logic'('1');
  --clock_crossing_0_m1_continuerequest continued request, which is an e_assign
  clock_crossing_0_m1_continuerequest <= std_logic'('1');
  internal_clock_crossing_0_m1_qualified_request_button_pio_s1 <= internal_clock_crossing_0_m1_requests_button_pio_s1 AND NOT ((clock_crossing_0_m1_read AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(clock_crossing_0_m1_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))))));
  --local readdatavalid clock_crossing_0_m1_read_data_valid_button_pio_s1, which is an e_mux
  clock_crossing_0_m1_read_data_valid_button_pio_s1 <= (internal_clock_crossing_0_m1_granted_button_pio_s1 AND clock_crossing_0_m1_read) AND NOT button_pio_s1_waits_for_read;
  --master is always granted when requested
  internal_clock_crossing_0_m1_granted_button_pio_s1 <= internal_clock_crossing_0_m1_qualified_request_button_pio_s1;
  --clock_crossing_0/m1 saved-grant button_pio/s1, which is an e_assign
  clock_crossing_0_m1_saved_grant_button_pio_s1 <= internal_clock_crossing_0_m1_requests_button_pio_s1;
  --allow new arb cycle for button_pio/s1, which is an e_assign
  button_pio_s1_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  button_pio_s1_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  button_pio_s1_master_qreq_vector <= std_logic'('1');
  --button_pio_s1_reset_n assignment, which is an e_assign
  button_pio_s1_reset_n <= reset_n;
  --button_pio_s1_firsttransfer first transaction, which is an e_assign
  button_pio_s1_firsttransfer <= A_WE_StdLogic((std_logic'(button_pio_s1_begins_xfer) = '1'), button_pio_s1_unreg_firsttransfer, button_pio_s1_reg_firsttransfer);
  --button_pio_s1_unreg_firsttransfer first transaction, which is an e_assign
  button_pio_s1_unreg_firsttransfer <= NOT ((button_pio_s1_slavearbiterlockenable AND button_pio_s1_any_continuerequest));
  --button_pio_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      button_pio_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(button_pio_s1_begins_xfer) = '1' then 
        button_pio_s1_reg_firsttransfer <= button_pio_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --button_pio_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  button_pio_s1_beginbursttransfer_internal <= button_pio_s1_begins_xfer;
  --button_pio_s1_address mux, which is an e_mux
  button_pio_s1_address <= clock_crossing_0_m1_nativeaddress (1 DOWNTO 0);
  --d1_button_pio_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_button_pio_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_button_pio_s1_end_xfer <= button_pio_s1_end_xfer;
    end if;

  end process;

  --button_pio_s1_waits_for_read in a cycle, which is an e_mux
  button_pio_s1_waits_for_read <= button_pio_s1_in_a_read_cycle AND button_pio_s1_begins_xfer;
  --button_pio_s1_in_a_read_cycle assignment, which is an e_assign
  button_pio_s1_in_a_read_cycle <= internal_clock_crossing_0_m1_granted_button_pio_s1 AND clock_crossing_0_m1_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= button_pio_s1_in_a_read_cycle;
  --button_pio_s1_waits_for_write in a cycle, which is an e_mux
  button_pio_s1_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(button_pio_s1_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --button_pio_s1_in_a_write_cycle assignment, which is an e_assign
  button_pio_s1_in_a_write_cycle <= internal_clock_crossing_0_m1_granted_button_pio_s1 AND clock_crossing_0_m1_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= button_pio_s1_in_a_write_cycle;
  wait_for_button_pio_s1_counter <= std_logic'('0');
  --vhdl renameroo for output signals
  clock_crossing_0_m1_granted_button_pio_s1 <= internal_clock_crossing_0_m1_granted_button_pio_s1;
  --vhdl renameroo for output signals
  clock_crossing_0_m1_qualified_request_button_pio_s1 <= internal_clock_crossing_0_m1_qualified_request_button_pio_s1;
  --vhdl renameroo for output signals
  clock_crossing_0_m1_requests_button_pio_s1 <= internal_clock_crossing_0_m1_requests_button_pio_s1;
--synthesis translate_off
    --button_pio/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity rdv_fifo_for_pcp_cpu_data_master_to_clock_crossing_0_s1_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC;
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity rdv_fifo_for_pcp_cpu_data_master_to_clock_crossing_0_s1_module;


architecture europa of rdv_fifo_for_pcp_cpu_data_master_to_clock_crossing_0_s1_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_10 :  STD_LOGIC;
                signal full_11 :  STD_LOGIC;
                signal full_12 :  STD_LOGIC;
                signal full_13 :  STD_LOGIC;
                signal full_14 :  STD_LOGIC;
                signal full_15 :  STD_LOGIC;
                signal full_16 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal full_3 :  STD_LOGIC;
                signal full_4 :  STD_LOGIC;
                signal full_5 :  STD_LOGIC;
                signal full_6 :  STD_LOGIC;
                signal full_7 :  STD_LOGIC;
                signal full_8 :  STD_LOGIC;
                signal full_9 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC;
                signal p10_full_10 :  STD_LOGIC;
                signal p10_stage_10 :  STD_LOGIC;
                signal p11_full_11 :  STD_LOGIC;
                signal p11_stage_11 :  STD_LOGIC;
                signal p12_full_12 :  STD_LOGIC;
                signal p12_stage_12 :  STD_LOGIC;
                signal p13_full_13 :  STD_LOGIC;
                signal p13_stage_13 :  STD_LOGIC;
                signal p14_full_14 :  STD_LOGIC;
                signal p14_stage_14 :  STD_LOGIC;
                signal p15_full_15 :  STD_LOGIC;
                signal p15_stage_15 :  STD_LOGIC;
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC;
                signal p2_full_2 :  STD_LOGIC;
                signal p2_stage_2 :  STD_LOGIC;
                signal p3_full_3 :  STD_LOGIC;
                signal p3_stage_3 :  STD_LOGIC;
                signal p4_full_4 :  STD_LOGIC;
                signal p4_stage_4 :  STD_LOGIC;
                signal p5_full_5 :  STD_LOGIC;
                signal p5_stage_5 :  STD_LOGIC;
                signal p6_full_6 :  STD_LOGIC;
                signal p6_stage_6 :  STD_LOGIC;
                signal p7_full_7 :  STD_LOGIC;
                signal p7_stage_7 :  STD_LOGIC;
                signal p8_full_8 :  STD_LOGIC;
                signal p8_stage_8 :  STD_LOGIC;
                signal p9_full_9 :  STD_LOGIC;
                signal p9_stage_9 :  STD_LOGIC;
                signal stage_0 :  STD_LOGIC;
                signal stage_1 :  STD_LOGIC;
                signal stage_10 :  STD_LOGIC;
                signal stage_11 :  STD_LOGIC;
                signal stage_12 :  STD_LOGIC;
                signal stage_13 :  STD_LOGIC;
                signal stage_14 :  STD_LOGIC;
                signal stage_15 :  STD_LOGIC;
                signal stage_2 :  STD_LOGIC;
                signal stage_3 :  STD_LOGIC;
                signal stage_4 :  STD_LOGIC;
                signal stage_5 :  STD_LOGIC;
                signal stage_6 :  STD_LOGIC;
                signal stage_7 :  STD_LOGIC;
                signal stage_8 :  STD_LOGIC;
                signal stage_9 :  STD_LOGIC;
                signal updated_one_count :  STD_LOGIC_VECTOR (5 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_15;
  empty <= NOT(full_0);
  full_16 <= std_logic'('0');
  --data_15, which is an e_mux
  p15_stage_15 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_16 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_15, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_15 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_15))))) = '1' then 
        if std_logic'(((sync_reset AND full_15) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_16))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_15 <= std_logic'('0');
        else
          stage_15 <= p15_stage_15;
        end if;
      end if;
    end if;

  end process;

  --control_15, which is an e_mux
  p15_full_15 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_14))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_15, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_15 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_15 <= std_logic'('0');
        else
          full_15 <= p15_full_15;
        end if;
      end if;
    end if;

  end process;

  --data_14, which is an e_mux
  p14_stage_14 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_15 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_15);
  --data_reg_14, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_14 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_14))))) = '1' then 
        if std_logic'(((sync_reset AND full_14) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_15))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_14 <= std_logic'('0');
        else
          stage_14 <= p14_stage_14;
        end if;
      end if;
    end if;

  end process;

  --control_14, which is an e_mux
  p14_full_14 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_13, full_15);
  --control_reg_14, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_14 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_14 <= std_logic'('0');
        else
          full_14 <= p14_full_14;
        end if;
      end if;
    end if;

  end process;

  --data_13, which is an e_mux
  p13_stage_13 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_14 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_14);
  --data_reg_13, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_13 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_13))))) = '1' then 
        if std_logic'(((sync_reset AND full_13) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_14))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_13 <= std_logic'('0');
        else
          stage_13 <= p13_stage_13;
        end if;
      end if;
    end if;

  end process;

  --control_13, which is an e_mux
  p13_full_13 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_12, full_14);
  --control_reg_13, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_13 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_13 <= std_logic'('0');
        else
          full_13 <= p13_full_13;
        end if;
      end if;
    end if;

  end process;

  --data_12, which is an e_mux
  p12_stage_12 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_13 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_13);
  --data_reg_12, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_12 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_12))))) = '1' then 
        if std_logic'(((sync_reset AND full_12) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_13))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_12 <= std_logic'('0');
        else
          stage_12 <= p12_stage_12;
        end if;
      end if;
    end if;

  end process;

  --control_12, which is an e_mux
  p12_full_12 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_11, full_13);
  --control_reg_12, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_12 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_12 <= std_logic'('0');
        else
          full_12 <= p12_full_12;
        end if;
      end if;
    end if;

  end process;

  --data_11, which is an e_mux
  p11_stage_11 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_12 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_12);
  --data_reg_11, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_11 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_11))))) = '1' then 
        if std_logic'(((sync_reset AND full_11) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_12))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_11 <= std_logic'('0');
        else
          stage_11 <= p11_stage_11;
        end if;
      end if;
    end if;

  end process;

  --control_11, which is an e_mux
  p11_full_11 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_10, full_12);
  --control_reg_11, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_11 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_11 <= std_logic'('0');
        else
          full_11 <= p11_full_11;
        end if;
      end if;
    end if;

  end process;

  --data_10, which is an e_mux
  p10_stage_10 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_11 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_11);
  --data_reg_10, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_10 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_10))))) = '1' then 
        if std_logic'(((sync_reset AND full_10) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_11))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_10 <= std_logic'('0');
        else
          stage_10 <= p10_stage_10;
        end if;
      end if;
    end if;

  end process;

  --control_10, which is an e_mux
  p10_full_10 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_9, full_11);
  --control_reg_10, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_10 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_10 <= std_logic'('0');
        else
          full_10 <= p10_full_10;
        end if;
      end if;
    end if;

  end process;

  --data_9, which is an e_mux
  p9_stage_9 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_10 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_10);
  --data_reg_9, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_9 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_9))))) = '1' then 
        if std_logic'(((sync_reset AND full_9) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_10))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_9 <= std_logic'('0');
        else
          stage_9 <= p9_stage_9;
        end if;
      end if;
    end if;

  end process;

  --control_9, which is an e_mux
  p9_full_9 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_8, full_10);
  --control_reg_9, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_9 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_9 <= std_logic'('0');
        else
          full_9 <= p9_full_9;
        end if;
      end if;
    end if;

  end process;

  --data_8, which is an e_mux
  p8_stage_8 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_9 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_9);
  --data_reg_8, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_8 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_8))))) = '1' then 
        if std_logic'(((sync_reset AND full_8) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_9))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_8 <= std_logic'('0');
        else
          stage_8 <= p8_stage_8;
        end if;
      end if;
    end if;

  end process;

  --control_8, which is an e_mux
  p8_full_8 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_7, full_9);
  --control_reg_8, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_8 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_8 <= std_logic'('0');
        else
          full_8 <= p8_full_8;
        end if;
      end if;
    end if;

  end process;

  --data_7, which is an e_mux
  p7_stage_7 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_8 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_8);
  --data_reg_7, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_7 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_7))))) = '1' then 
        if std_logic'(((sync_reset AND full_7) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_8))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_7 <= std_logic'('0');
        else
          stage_7 <= p7_stage_7;
        end if;
      end if;
    end if;

  end process;

  --control_7, which is an e_mux
  p7_full_7 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_6, full_8);
  --control_reg_7, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_7 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_7 <= std_logic'('0');
        else
          full_7 <= p7_full_7;
        end if;
      end if;
    end if;

  end process;

  --data_6, which is an e_mux
  p6_stage_6 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_7 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_7);
  --data_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_6 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_6))))) = '1' then 
        if std_logic'(((sync_reset AND full_6) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_7))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_6 <= std_logic'('0');
        else
          stage_6 <= p6_stage_6;
        end if;
      end if;
    end if;

  end process;

  --control_6, which is an e_mux
  p6_full_6 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_5, full_7);
  --control_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_6 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_6 <= std_logic'('0');
        else
          full_6 <= p6_full_6;
        end if;
      end if;
    end if;

  end process;

  --data_5, which is an e_mux
  p5_stage_5 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_6 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_6);
  --data_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_5))))) = '1' then 
        if std_logic'(((sync_reset AND full_5) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_6))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_5 <= std_logic'('0');
        else
          stage_5 <= p5_stage_5;
        end if;
      end if;
    end if;

  end process;

  --control_5, which is an e_mux
  p5_full_5 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_4, full_6);
  --control_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_5 <= std_logic'('0');
        else
          full_5 <= p5_full_5;
        end if;
      end if;
    end if;

  end process;

  --data_4, which is an e_mux
  p4_stage_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_5 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_5);
  --data_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_4))))) = '1' then 
        if std_logic'(((sync_reset AND full_4) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_5))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_4 <= std_logic'('0');
        else
          stage_4 <= p4_stage_4;
        end if;
      end if;
    end if;

  end process;

  --control_4, which is an e_mux
  p4_full_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_3, full_5);
  --control_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_4 <= std_logic'('0');
        else
          full_4 <= p4_full_4;
        end if;
      end if;
    end if;

  end process;

  --data_3, which is an e_mux
  p3_stage_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_4 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_4);
  --data_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_3))))) = '1' then 
        if std_logic'(((sync_reset AND full_3) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_4))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_3 <= std_logic'('0');
        else
          stage_3 <= p3_stage_3;
        end if;
      end if;
    end if;

  end process;

  --control_3, which is an e_mux
  p3_full_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_2, full_4);
  --control_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_3 <= std_logic'('0');
        else
          full_3 <= p3_full_3;
        end if;
      end if;
    end if;

  end process;

  --data_2, which is an e_mux
  p2_stage_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_3 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_3);
  --data_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_2))))) = '1' then 
        if std_logic'(((sync_reset AND full_2) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_3))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_2 <= std_logic'('0');
        else
          stage_2 <= p2_stage_2;
        end if;
      end if;
    end if;

  end process;

  --control_2, which is an e_mux
  p2_full_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_1, full_3);
  --control_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_2 <= std_logic'('0');
        else
          full_2 <= p2_full_2;
        end if;
      end if;
    end if;

  end process;

  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_2);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic'('0');
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_0, full_2);
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic'('0');
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 6);
  one_count_minus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 6);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("00000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("00000") & (A_TOSTDLOGICVECTOR(data_in))), A_WE_StdLogicVector((std_logic'(((((read AND (data_in)) AND write) AND (stage_0)))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (data_in)))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (stage_0)))) = '1'), one_count_minus_one, how_many_ones))))))), 6);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity clock_crossing_0_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal clock_crossing_0_s1_endofpacket : IN STD_LOGIC;
                 signal clock_crossing_0_s1_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal clock_crossing_0_s1_readdatavalid : IN STD_LOGIC;
                 signal clock_crossing_0_s1_waitrequest : IN STD_LOGIC;
                 signal pcp_cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (25 DOWNTO 0);
                 signal pcp_cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal pcp_cpu_data_master_read : IN STD_LOGIC;
                 signal pcp_cpu_data_master_waitrequest : IN STD_LOGIC;
                 signal pcp_cpu_data_master_write : IN STD_LOGIC;
                 signal pcp_cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal clock_crossing_0_s1_address : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
                 signal clock_crossing_0_s1_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal clock_crossing_0_s1_endofpacket_from_sa : OUT STD_LOGIC;
                 signal clock_crossing_0_s1_nativeaddress : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
                 signal clock_crossing_0_s1_read : OUT STD_LOGIC;
                 signal clock_crossing_0_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal clock_crossing_0_s1_reset_n : OUT STD_LOGIC;
                 signal clock_crossing_0_s1_waitrequest_from_sa : OUT STD_LOGIC;
                 signal clock_crossing_0_s1_write : OUT STD_LOGIC;
                 signal clock_crossing_0_s1_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal d1_clock_crossing_0_s1_end_xfer : OUT STD_LOGIC;
                 signal pcp_cpu_data_master_granted_clock_crossing_0_s1 : OUT STD_LOGIC;
                 signal pcp_cpu_data_master_qualified_request_clock_crossing_0_s1 : OUT STD_LOGIC;
                 signal pcp_cpu_data_master_read_data_valid_clock_crossing_0_s1 : OUT STD_LOGIC;
                 signal pcp_cpu_data_master_read_data_valid_clock_crossing_0_s1_shift_register : OUT STD_LOGIC;
                 signal pcp_cpu_data_master_requests_clock_crossing_0_s1 : OUT STD_LOGIC
              );
end entity clock_crossing_0_s1_arbitrator;


architecture europa of clock_crossing_0_s1_arbitrator is
component rdv_fifo_for_pcp_cpu_data_master_to_clock_crossing_0_s1_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC;
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component rdv_fifo_for_pcp_cpu_data_master_to_clock_crossing_0_s1_module;

                signal clock_crossing_0_s1_allgrants :  STD_LOGIC;
                signal clock_crossing_0_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal clock_crossing_0_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal clock_crossing_0_s1_any_continuerequest :  STD_LOGIC;
                signal clock_crossing_0_s1_arb_counter_enable :  STD_LOGIC;
                signal clock_crossing_0_s1_arb_share_counter :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal clock_crossing_0_s1_arb_share_counter_next_value :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal clock_crossing_0_s1_arb_share_set_values :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal clock_crossing_0_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal clock_crossing_0_s1_begins_xfer :  STD_LOGIC;
                signal clock_crossing_0_s1_end_xfer :  STD_LOGIC;
                signal clock_crossing_0_s1_firsttransfer :  STD_LOGIC;
                signal clock_crossing_0_s1_grant_vector :  STD_LOGIC;
                signal clock_crossing_0_s1_in_a_read_cycle :  STD_LOGIC;
                signal clock_crossing_0_s1_in_a_write_cycle :  STD_LOGIC;
                signal clock_crossing_0_s1_master_qreq_vector :  STD_LOGIC;
                signal clock_crossing_0_s1_move_on_to_next_transaction :  STD_LOGIC;
                signal clock_crossing_0_s1_non_bursting_master_requests :  STD_LOGIC;
                signal clock_crossing_0_s1_readdatavalid_from_sa :  STD_LOGIC;
                signal clock_crossing_0_s1_reg_firsttransfer :  STD_LOGIC;
                signal clock_crossing_0_s1_slavearbiterlockenable :  STD_LOGIC;
                signal clock_crossing_0_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal clock_crossing_0_s1_unreg_firsttransfer :  STD_LOGIC;
                signal clock_crossing_0_s1_waits_for_read :  STD_LOGIC;
                signal clock_crossing_0_s1_waits_for_write :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_clock_crossing_0_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_clock_crossing_0_s1_waitrequest_from_sa :  STD_LOGIC;
                signal internal_pcp_cpu_data_master_granted_clock_crossing_0_s1 :  STD_LOGIC;
                signal internal_pcp_cpu_data_master_qualified_request_clock_crossing_0_s1 :  STD_LOGIC;
                signal internal_pcp_cpu_data_master_read_data_valid_clock_crossing_0_s1_shift_register :  STD_LOGIC;
                signal internal_pcp_cpu_data_master_requests_clock_crossing_0_s1 :  STD_LOGIC;
                signal module_input :  STD_LOGIC;
                signal module_input1 :  STD_LOGIC;
                signal module_input2 :  STD_LOGIC;
                signal pcp_cpu_data_master_arbiterlock :  STD_LOGIC;
                signal pcp_cpu_data_master_arbiterlock2 :  STD_LOGIC;
                signal pcp_cpu_data_master_continuerequest :  STD_LOGIC;
                signal pcp_cpu_data_master_rdv_fifo_empty_clock_crossing_0_s1 :  STD_LOGIC;
                signal pcp_cpu_data_master_rdv_fifo_output_from_clock_crossing_0_s1 :  STD_LOGIC;
                signal pcp_cpu_data_master_saved_grant_clock_crossing_0_s1 :  STD_LOGIC;
                signal shifted_address_to_clock_crossing_0_s1_from_pcp_cpu_data_master :  STD_LOGIC_VECTOR (25 DOWNTO 0);
                signal wait_for_clock_crossing_0_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT clock_crossing_0_s1_end_xfer;
    end if;

  end process;

  clock_crossing_0_s1_begins_xfer <= NOT d1_reasons_to_wait AND (internal_pcp_cpu_data_master_qualified_request_clock_crossing_0_s1);
  --assign clock_crossing_0_s1_readdata_from_sa = clock_crossing_0_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  clock_crossing_0_s1_readdata_from_sa <= clock_crossing_0_s1_readdata;
  internal_pcp_cpu_data_master_requests_clock_crossing_0_s1 <= to_std_logic(((Std_Logic_Vector'(pcp_cpu_data_master_address_to_slave(25 DOWNTO 7) & std_logic_vector'("0000000")) = std_logic_vector'("01000000000000000000000000")))) AND ((pcp_cpu_data_master_read OR pcp_cpu_data_master_write));
  --assign clock_crossing_0_s1_waitrequest_from_sa = clock_crossing_0_s1_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_clock_crossing_0_s1_waitrequest_from_sa <= clock_crossing_0_s1_waitrequest;
  --assign clock_crossing_0_s1_readdatavalid_from_sa = clock_crossing_0_s1_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  clock_crossing_0_s1_readdatavalid_from_sa <= clock_crossing_0_s1_readdatavalid;
  --clock_crossing_0_s1_arb_share_counter set values, which is an e_mux
  clock_crossing_0_s1_arb_share_set_values <= std_logic_vector'("01");
  --clock_crossing_0_s1_non_bursting_master_requests mux, which is an e_mux
  clock_crossing_0_s1_non_bursting_master_requests <= internal_pcp_cpu_data_master_requests_clock_crossing_0_s1;
  --clock_crossing_0_s1_any_bursting_master_saved_grant mux, which is an e_mux
  clock_crossing_0_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --clock_crossing_0_s1_arb_share_counter_next_value assignment, which is an e_assign
  clock_crossing_0_s1_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(clock_crossing_0_s1_firsttransfer) = '1'), (((std_logic_vector'("0000000000000000000000000000000") & (clock_crossing_0_s1_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(clock_crossing_0_s1_arb_share_counter)) = '1'), (((std_logic_vector'("0000000000000000000000000000000") & (clock_crossing_0_s1_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 2);
  --clock_crossing_0_s1_allgrants all slave grants, which is an e_mux
  clock_crossing_0_s1_allgrants <= clock_crossing_0_s1_grant_vector;
  --clock_crossing_0_s1_end_xfer assignment, which is an e_assign
  clock_crossing_0_s1_end_xfer <= NOT ((clock_crossing_0_s1_waits_for_read OR clock_crossing_0_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_clock_crossing_0_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_clock_crossing_0_s1 <= clock_crossing_0_s1_end_xfer AND (((NOT clock_crossing_0_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --clock_crossing_0_s1_arb_share_counter arbitration counter enable, which is an e_assign
  clock_crossing_0_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_clock_crossing_0_s1 AND clock_crossing_0_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_clock_crossing_0_s1 AND NOT clock_crossing_0_s1_non_bursting_master_requests));
  --clock_crossing_0_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      clock_crossing_0_s1_arb_share_counter <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      if std_logic'(clock_crossing_0_s1_arb_counter_enable) = '1' then 
        clock_crossing_0_s1_arb_share_counter <= clock_crossing_0_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --clock_crossing_0_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      clock_crossing_0_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clock_crossing_0_s1_master_qreq_vector AND end_xfer_arb_share_counter_term_clock_crossing_0_s1)) OR ((end_xfer_arb_share_counter_term_clock_crossing_0_s1 AND NOT clock_crossing_0_s1_non_bursting_master_requests)))) = '1' then 
        clock_crossing_0_s1_slavearbiterlockenable <= or_reduce(clock_crossing_0_s1_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --pcp_cpu/data_master clock_crossing_0/s1 arbiterlock, which is an e_assign
  pcp_cpu_data_master_arbiterlock <= clock_crossing_0_s1_slavearbiterlockenable AND pcp_cpu_data_master_continuerequest;
  --clock_crossing_0_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  clock_crossing_0_s1_slavearbiterlockenable2 <= or_reduce(clock_crossing_0_s1_arb_share_counter_next_value);
  --pcp_cpu/data_master clock_crossing_0/s1 arbiterlock2, which is an e_assign
  pcp_cpu_data_master_arbiterlock2 <= clock_crossing_0_s1_slavearbiterlockenable2 AND pcp_cpu_data_master_continuerequest;
  --clock_crossing_0_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  clock_crossing_0_s1_any_continuerequest <= std_logic'('1');
  --pcp_cpu_data_master_continuerequest continued request, which is an e_assign
  pcp_cpu_data_master_continuerequest <= std_logic'('1');
  internal_pcp_cpu_data_master_qualified_request_clock_crossing_0_s1 <= internal_pcp_cpu_data_master_requests_clock_crossing_0_s1 AND NOT ((((pcp_cpu_data_master_read AND ((NOT pcp_cpu_data_master_waitrequest OR (internal_pcp_cpu_data_master_read_data_valid_clock_crossing_0_s1_shift_register))))) OR (((NOT pcp_cpu_data_master_waitrequest) AND pcp_cpu_data_master_write))));
  --unique name for clock_crossing_0_s1_move_on_to_next_transaction, which is an e_assign
  clock_crossing_0_s1_move_on_to_next_transaction <= clock_crossing_0_s1_readdatavalid_from_sa;
  --rdv_fifo_for_pcp_cpu_data_master_to_clock_crossing_0_s1, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_pcp_cpu_data_master_to_clock_crossing_0_s1 : rdv_fifo_for_pcp_cpu_data_master_to_clock_crossing_0_s1_module
    port map(
      data_out => pcp_cpu_data_master_rdv_fifo_output_from_clock_crossing_0_s1,
      empty => open,
      fifo_contains_ones_n => pcp_cpu_data_master_rdv_fifo_empty_clock_crossing_0_s1,
      full => open,
      clear_fifo => module_input,
      clk => clk,
      data_in => internal_pcp_cpu_data_master_granted_clock_crossing_0_s1,
      read => clock_crossing_0_s1_move_on_to_next_transaction,
      reset_n => reset_n,
      sync_reset => module_input1,
      write => module_input2
    );

  module_input <= std_logic'('0');
  module_input1 <= std_logic'('0');
  module_input2 <= in_a_read_cycle AND NOT clock_crossing_0_s1_waits_for_read;

  internal_pcp_cpu_data_master_read_data_valid_clock_crossing_0_s1_shift_register <= NOT pcp_cpu_data_master_rdv_fifo_empty_clock_crossing_0_s1;
  --local readdatavalid pcp_cpu_data_master_read_data_valid_clock_crossing_0_s1, which is an e_mux
  pcp_cpu_data_master_read_data_valid_clock_crossing_0_s1 <= clock_crossing_0_s1_readdatavalid_from_sa;
  --clock_crossing_0_s1_writedata mux, which is an e_mux
  clock_crossing_0_s1_writedata <= pcp_cpu_data_master_writedata;
  --assign clock_crossing_0_s1_endofpacket_from_sa = clock_crossing_0_s1_endofpacket so that symbol knows where to group signals which may go to master only, which is an e_assign
  clock_crossing_0_s1_endofpacket_from_sa <= clock_crossing_0_s1_endofpacket;
  --master is always granted when requested
  internal_pcp_cpu_data_master_granted_clock_crossing_0_s1 <= internal_pcp_cpu_data_master_qualified_request_clock_crossing_0_s1;
  --pcp_cpu/data_master saved-grant clock_crossing_0/s1, which is an e_assign
  pcp_cpu_data_master_saved_grant_clock_crossing_0_s1 <= internal_pcp_cpu_data_master_requests_clock_crossing_0_s1;
  --allow new arb cycle for clock_crossing_0/s1, which is an e_assign
  clock_crossing_0_s1_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  clock_crossing_0_s1_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  clock_crossing_0_s1_master_qreq_vector <= std_logic'('1');
  --clock_crossing_0_s1_reset_n assignment, which is an e_assign
  clock_crossing_0_s1_reset_n <= reset_n;
  --clock_crossing_0_s1_firsttransfer first transaction, which is an e_assign
  clock_crossing_0_s1_firsttransfer <= A_WE_StdLogic((std_logic'(clock_crossing_0_s1_begins_xfer) = '1'), clock_crossing_0_s1_unreg_firsttransfer, clock_crossing_0_s1_reg_firsttransfer);
  --clock_crossing_0_s1_unreg_firsttransfer first transaction, which is an e_assign
  clock_crossing_0_s1_unreg_firsttransfer <= NOT ((clock_crossing_0_s1_slavearbiterlockenable AND clock_crossing_0_s1_any_continuerequest));
  --clock_crossing_0_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      clock_crossing_0_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(clock_crossing_0_s1_begins_xfer) = '1' then 
        clock_crossing_0_s1_reg_firsttransfer <= clock_crossing_0_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --clock_crossing_0_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  clock_crossing_0_s1_beginbursttransfer_internal <= clock_crossing_0_s1_begins_xfer;
  --clock_crossing_0_s1_read assignment, which is an e_mux
  clock_crossing_0_s1_read <= internal_pcp_cpu_data_master_granted_clock_crossing_0_s1 AND pcp_cpu_data_master_read;
  --clock_crossing_0_s1_write assignment, which is an e_mux
  clock_crossing_0_s1_write <= internal_pcp_cpu_data_master_granted_clock_crossing_0_s1 AND pcp_cpu_data_master_write;
  shifted_address_to_clock_crossing_0_s1_from_pcp_cpu_data_master <= pcp_cpu_data_master_address_to_slave;
  --clock_crossing_0_s1_address mux, which is an e_mux
  clock_crossing_0_s1_address <= A_EXT (A_SRL(shifted_address_to_clock_crossing_0_s1_from_pcp_cpu_data_master,std_logic_vector'("00000000000000000000000000000010")), 5);
  --slaveid clock_crossing_0_s1_nativeaddress nativeaddress mux, which is an e_mux
  clock_crossing_0_s1_nativeaddress <= A_EXT (A_SRL(pcp_cpu_data_master_address_to_slave,std_logic_vector'("00000000000000000000000000000010")), 5);
  --d1_clock_crossing_0_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_clock_crossing_0_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_clock_crossing_0_s1_end_xfer <= clock_crossing_0_s1_end_xfer;
    end if;

  end process;

  --clock_crossing_0_s1_waits_for_read in a cycle, which is an e_mux
  clock_crossing_0_s1_waits_for_read <= clock_crossing_0_s1_in_a_read_cycle AND internal_clock_crossing_0_s1_waitrequest_from_sa;
  --clock_crossing_0_s1_in_a_read_cycle assignment, which is an e_assign
  clock_crossing_0_s1_in_a_read_cycle <= internal_pcp_cpu_data_master_granted_clock_crossing_0_s1 AND pcp_cpu_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= clock_crossing_0_s1_in_a_read_cycle;
  --clock_crossing_0_s1_waits_for_write in a cycle, which is an e_mux
  clock_crossing_0_s1_waits_for_write <= clock_crossing_0_s1_in_a_write_cycle AND internal_clock_crossing_0_s1_waitrequest_from_sa;
  --clock_crossing_0_s1_in_a_write_cycle assignment, which is an e_assign
  clock_crossing_0_s1_in_a_write_cycle <= internal_pcp_cpu_data_master_granted_clock_crossing_0_s1 AND pcp_cpu_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= clock_crossing_0_s1_in_a_write_cycle;
  wait_for_clock_crossing_0_s1_counter <= std_logic'('0');
  --clock_crossing_0_s1_byteenable byte enable port mux, which is an e_mux
  clock_crossing_0_s1_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_pcp_cpu_data_master_granted_clock_crossing_0_s1)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (pcp_cpu_data_master_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))), 4);
  --vhdl renameroo for output signals
  clock_crossing_0_s1_waitrequest_from_sa <= internal_clock_crossing_0_s1_waitrequest_from_sa;
  --vhdl renameroo for output signals
  pcp_cpu_data_master_granted_clock_crossing_0_s1 <= internal_pcp_cpu_data_master_granted_clock_crossing_0_s1;
  --vhdl renameroo for output signals
  pcp_cpu_data_master_qualified_request_clock_crossing_0_s1 <= internal_pcp_cpu_data_master_qualified_request_clock_crossing_0_s1;
  --vhdl renameroo for output signals
  pcp_cpu_data_master_read_data_valid_clock_crossing_0_s1_shift_register <= internal_pcp_cpu_data_master_read_data_valid_clock_crossing_0_s1_shift_register;
  --vhdl renameroo for output signals
  pcp_cpu_data_master_requests_clock_crossing_0_s1 <= internal_pcp_cpu_data_master_requests_clock_crossing_0_s1;
--synthesis translate_off
    --clock_crossing_0/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity clock_crossing_0_m1_arbitrator is 
        port (
              -- inputs:
                 signal button_pio_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal clk : IN STD_LOGIC;
                 signal clock_crossing_0_m1_address : IN STD_LOGIC_VECTOR (6 DOWNTO 0);
                 signal clock_crossing_0_m1_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal clock_crossing_0_m1_granted_button_pio_s1 : IN STD_LOGIC;
                 signal clock_crossing_0_m1_granted_irq_gen_s1 : IN STD_LOGIC;
                 signal clock_crossing_0_m1_granted_status_led_pio_s1 : IN STD_LOGIC;
                 signal clock_crossing_0_m1_granted_sysid_control_slave : IN STD_LOGIC;
                 signal clock_crossing_0_m1_granted_system_timer_s1 : IN STD_LOGIC;
                 signal clock_crossing_0_m1_qualified_request_button_pio_s1 : IN STD_LOGIC;
                 signal clock_crossing_0_m1_qualified_request_irq_gen_s1 : IN STD_LOGIC;
                 signal clock_crossing_0_m1_qualified_request_status_led_pio_s1 : IN STD_LOGIC;
                 signal clock_crossing_0_m1_qualified_request_sysid_control_slave : IN STD_LOGIC;
                 signal clock_crossing_0_m1_qualified_request_system_timer_s1 : IN STD_LOGIC;
                 signal clock_crossing_0_m1_read : IN STD_LOGIC;
                 signal clock_crossing_0_m1_read_data_valid_button_pio_s1 : IN STD_LOGIC;
                 signal clock_crossing_0_m1_read_data_valid_irq_gen_s1 : IN STD_LOGIC;
                 signal clock_crossing_0_m1_read_data_valid_status_led_pio_s1 : IN STD_LOGIC;
                 signal clock_crossing_0_m1_read_data_valid_sysid_control_slave : IN STD_LOGIC;
                 signal clock_crossing_0_m1_read_data_valid_system_timer_s1 : IN STD_LOGIC;
                 signal clock_crossing_0_m1_requests_button_pio_s1 : IN STD_LOGIC;
                 signal clock_crossing_0_m1_requests_irq_gen_s1 : IN STD_LOGIC;
                 signal clock_crossing_0_m1_requests_status_led_pio_s1 : IN STD_LOGIC;
                 signal clock_crossing_0_m1_requests_sysid_control_slave : IN STD_LOGIC;
                 signal clock_crossing_0_m1_requests_system_timer_s1 : IN STD_LOGIC;
                 signal clock_crossing_0_m1_write : IN STD_LOGIC;
                 signal clock_crossing_0_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal d1_button_pio_s1_end_xfer : IN STD_LOGIC;
                 signal d1_irq_gen_s1_end_xfer : IN STD_LOGIC;
                 signal d1_status_led_pio_s1_end_xfer : IN STD_LOGIC;
                 signal d1_sysid_control_slave_end_xfer : IN STD_LOGIC;
                 signal d1_system_timer_s1_end_xfer : IN STD_LOGIC;
                 signal irq_gen_s1_readdata_from_sa : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal status_led_pio_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal sysid_control_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal system_timer_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

              -- outputs:
                 signal clock_crossing_0_m1_address_to_slave : OUT STD_LOGIC_VECTOR (6 DOWNTO 0);
                 signal clock_crossing_0_m1_latency_counter : OUT STD_LOGIC;
                 signal clock_crossing_0_m1_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal clock_crossing_0_m1_readdatavalid : OUT STD_LOGIC;
                 signal clock_crossing_0_m1_reset_n : OUT STD_LOGIC;
                 signal clock_crossing_0_m1_waitrequest : OUT STD_LOGIC
              );
end entity clock_crossing_0_m1_arbitrator;


architecture europa of clock_crossing_0_m1_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal clock_crossing_0_m1_address_last_time :  STD_LOGIC_VECTOR (6 DOWNTO 0);
                signal clock_crossing_0_m1_byteenable_last_time :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal clock_crossing_0_m1_is_granted_some_slave :  STD_LOGIC;
                signal clock_crossing_0_m1_read_but_no_slave_selected :  STD_LOGIC;
                signal clock_crossing_0_m1_read_last_time :  STD_LOGIC;
                signal clock_crossing_0_m1_run :  STD_LOGIC;
                signal clock_crossing_0_m1_write_last_time :  STD_LOGIC;
                signal clock_crossing_0_m1_writedata_last_time :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal internal_clock_crossing_0_m1_address_to_slave :  STD_LOGIC_VECTOR (6 DOWNTO 0);
                signal internal_clock_crossing_0_m1_latency_counter :  STD_LOGIC;
                signal internal_clock_crossing_0_m1_waitrequest :  STD_LOGIC;
                signal latency_load_value :  STD_LOGIC;
                signal p1_clock_crossing_0_m1_latency_counter :  STD_LOGIC;
                signal pre_flush_clock_crossing_0_m1_readdatavalid :  STD_LOGIC;
                signal r_0 :  STD_LOGIC;
                signal r_2 :  STD_LOGIC;

begin

  --r_0 master_run cascaded wait assignment, which is an e_assign
  r_0 <= Vector_To_Std_Logic((((((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((clock_crossing_0_m1_qualified_request_button_pio_s1 OR NOT clock_crossing_0_m1_requests_button_pio_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT clock_crossing_0_m1_qualified_request_button_pio_s1 OR NOT clock_crossing_0_m1_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT d1_button_pio_s1_end_xfer)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(clock_crossing_0_m1_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT clock_crossing_0_m1_qualified_request_button_pio_s1 OR NOT clock_crossing_0_m1_write)))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(clock_crossing_0_m1_write)))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((clock_crossing_0_m1_qualified_request_irq_gen_s1 OR NOT clock_crossing_0_m1_requests_irq_gen_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT clock_crossing_0_m1_qualified_request_irq_gen_s1 OR NOT clock_crossing_0_m1_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT d1_irq_gen_s1_end_xfer)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(clock_crossing_0_m1_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT clock_crossing_0_m1_qualified_request_irq_gen_s1 OR NOT clock_crossing_0_m1_write)))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(clock_crossing_0_m1_write)))))))));
  --cascaded wait assignment, which is an e_assign
  clock_crossing_0_m1_run <= r_0 AND r_2;
  --r_2 master_run cascaded wait assignment, which is an e_assign
  r_2 <= Vector_To_Std_Logic(((((((((((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((clock_crossing_0_m1_qualified_request_status_led_pio_s1 OR NOT clock_crossing_0_m1_requests_status_led_pio_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT clock_crossing_0_m1_qualified_request_status_led_pio_s1 OR NOT clock_crossing_0_m1_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT d1_status_led_pio_s1_end_xfer)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(clock_crossing_0_m1_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT clock_crossing_0_m1_qualified_request_status_led_pio_s1 OR NOT clock_crossing_0_m1_write)))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(clock_crossing_0_m1_write)))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((clock_crossing_0_m1_qualified_request_sysid_control_slave OR NOT clock_crossing_0_m1_requests_sysid_control_slave)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((clock_crossing_0_m1_granted_sysid_control_slave OR NOT clock_crossing_0_m1_qualified_request_sysid_control_slave)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT clock_crossing_0_m1_qualified_request_sysid_control_slave OR NOT clock_crossing_0_m1_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT d1_sysid_control_slave_end_xfer)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(clock_crossing_0_m1_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT clock_crossing_0_m1_qualified_request_sysid_control_slave OR NOT clock_crossing_0_m1_write)))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(clock_crossing_0_m1_write)))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((clock_crossing_0_m1_qualified_request_system_timer_s1 OR NOT clock_crossing_0_m1_requests_system_timer_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT clock_crossing_0_m1_qualified_request_system_timer_s1 OR NOT clock_crossing_0_m1_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT d1_system_timer_s1_end_xfer)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(clock_crossing_0_m1_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT clock_crossing_0_m1_qualified_request_system_timer_s1 OR NOT clock_crossing_0_m1_write)))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(clock_crossing_0_m1_write)))))))));
  --optimize select-logic by passing only those address bits which matter.
  internal_clock_crossing_0_m1_address_to_slave <= clock_crossing_0_m1_address(6 DOWNTO 0);
  --clock_crossing_0_m1_read_but_no_slave_selected assignment, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      clock_crossing_0_m1_read_but_no_slave_selected <= std_logic'('0');
    elsif clk'event and clk = '1' then
      clock_crossing_0_m1_read_but_no_slave_selected <= (clock_crossing_0_m1_read AND clock_crossing_0_m1_run) AND NOT clock_crossing_0_m1_is_granted_some_slave;
    end if;

  end process;

  --some slave is getting selected, which is an e_mux
  clock_crossing_0_m1_is_granted_some_slave <= (((clock_crossing_0_m1_granted_button_pio_s1 OR clock_crossing_0_m1_granted_irq_gen_s1) OR clock_crossing_0_m1_granted_status_led_pio_s1) OR clock_crossing_0_m1_granted_sysid_control_slave) OR clock_crossing_0_m1_granted_system_timer_s1;
  --latent slave read data valids which may be flushed, which is an e_mux
  pre_flush_clock_crossing_0_m1_readdatavalid <= std_logic'('0');
  --latent slave read data valid which is not flushed, which is an e_mux
  clock_crossing_0_m1_readdatavalid <= (((((((((((((clock_crossing_0_m1_read_but_no_slave_selected OR pre_flush_clock_crossing_0_m1_readdatavalid) OR clock_crossing_0_m1_read_data_valid_button_pio_s1) OR clock_crossing_0_m1_read_but_no_slave_selected) OR pre_flush_clock_crossing_0_m1_readdatavalid) OR clock_crossing_0_m1_read_data_valid_irq_gen_s1) OR clock_crossing_0_m1_read_but_no_slave_selected) OR pre_flush_clock_crossing_0_m1_readdatavalid) OR clock_crossing_0_m1_read_data_valid_status_led_pio_s1) OR clock_crossing_0_m1_read_but_no_slave_selected) OR pre_flush_clock_crossing_0_m1_readdatavalid) OR clock_crossing_0_m1_read_data_valid_sysid_control_slave) OR clock_crossing_0_m1_read_but_no_slave_selected) OR pre_flush_clock_crossing_0_m1_readdatavalid) OR clock_crossing_0_m1_read_data_valid_system_timer_s1;
  --clock_crossing_0/m1 readdata mux, which is an e_mux
  clock_crossing_0_m1_readdata <= (((((A_REP(NOT ((clock_crossing_0_m1_qualified_request_button_pio_s1 AND clock_crossing_0_m1_read)) , 32) OR (std_logic_vector'("000000000000000000000000") & (button_pio_s1_readdata_from_sa)))) AND ((A_REP(NOT ((clock_crossing_0_m1_qualified_request_irq_gen_s1 AND clock_crossing_0_m1_read)) , 32) OR (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(irq_gen_s1_readdata_from_sa)))))) AND ((A_REP(NOT ((clock_crossing_0_m1_qualified_request_status_led_pio_s1 AND clock_crossing_0_m1_read)) , 32) OR (std_logic_vector'("000000000000000000000000") & (status_led_pio_s1_readdata_from_sa))))) AND ((A_REP(NOT ((clock_crossing_0_m1_qualified_request_sysid_control_slave AND clock_crossing_0_m1_read)) , 32) OR sysid_control_slave_readdata_from_sa))) AND ((A_REP(NOT ((clock_crossing_0_m1_qualified_request_system_timer_s1 AND clock_crossing_0_m1_read)) , 32) OR (std_logic_vector'("0000000000000000") & (system_timer_s1_readdata_from_sa))));
  --actual waitrequest port, which is an e_assign
  internal_clock_crossing_0_m1_waitrequest <= NOT clock_crossing_0_m1_run;
  --latent max counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      internal_clock_crossing_0_m1_latency_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      internal_clock_crossing_0_m1_latency_counter <= p1_clock_crossing_0_m1_latency_counter;
    end if;

  end process;

  --latency counter load mux, which is an e_mux
  p1_clock_crossing_0_m1_latency_counter <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(((clock_crossing_0_m1_run AND clock_crossing_0_m1_read))) = '1'), (std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(latency_load_value))), A_WE_StdLogicVector((std_logic'((internal_clock_crossing_0_m1_latency_counter)) = '1'), ((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(internal_clock_crossing_0_m1_latency_counter))) - std_logic_vector'("000000000000000000000000000000001")), std_logic_vector'("000000000000000000000000000000000"))));
  --read latency load values, which is an e_mux
  latency_load_value <= std_logic'('0');
  --clock_crossing_0_m1_reset_n assignment, which is an e_assign
  clock_crossing_0_m1_reset_n <= reset_n;
  --vhdl renameroo for output signals
  clock_crossing_0_m1_address_to_slave <= internal_clock_crossing_0_m1_address_to_slave;
  --vhdl renameroo for output signals
  clock_crossing_0_m1_latency_counter <= internal_clock_crossing_0_m1_latency_counter;
  --vhdl renameroo for output signals
  clock_crossing_0_m1_waitrequest <= internal_clock_crossing_0_m1_waitrequest;
--synthesis translate_off
    --clock_crossing_0_m1_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        clock_crossing_0_m1_address_last_time <= std_logic_vector'("0000000");
      elsif clk'event and clk = '1' then
        clock_crossing_0_m1_address_last_time <= clock_crossing_0_m1_address;
      end if;

    end process;

    --clock_crossing_0/m1 waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_clock_crossing_0_m1_waitrequest AND ((clock_crossing_0_m1_read OR clock_crossing_0_m1_write));
      end if;

    end process;

    --clock_crossing_0_m1_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line4 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((clock_crossing_0_m1_address /= clock_crossing_0_m1_address_last_time))))) = '1' then 
          write(write_line4, now);
          write(write_line4, string'(": "));
          write(write_line4, string'("clock_crossing_0_m1_address did not heed wait!!!"));
          write(output, write_line4.all);
          deallocate (write_line4);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --clock_crossing_0_m1_byteenable check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        clock_crossing_0_m1_byteenable_last_time <= std_logic_vector'("0000");
      elsif clk'event and clk = '1' then
        clock_crossing_0_m1_byteenable_last_time <= clock_crossing_0_m1_byteenable;
      end if;

    end process;

    --clock_crossing_0_m1_byteenable matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line5 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((clock_crossing_0_m1_byteenable /= clock_crossing_0_m1_byteenable_last_time))))) = '1' then 
          write(write_line5, now);
          write(write_line5, string'(": "));
          write(write_line5, string'("clock_crossing_0_m1_byteenable did not heed wait!!!"));
          write(output, write_line5.all);
          deallocate (write_line5);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --clock_crossing_0_m1_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        clock_crossing_0_m1_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        clock_crossing_0_m1_read_last_time <= clock_crossing_0_m1_read;
      end if;

    end process;

    --clock_crossing_0_m1_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line6 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(clock_crossing_0_m1_read) /= std_logic'(clock_crossing_0_m1_read_last_time)))))) = '1' then 
          write(write_line6, now);
          write(write_line6, string'(": "));
          write(write_line6, string'("clock_crossing_0_m1_read did not heed wait!!!"));
          write(output, write_line6.all);
          deallocate (write_line6);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --clock_crossing_0_m1_write check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        clock_crossing_0_m1_write_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        clock_crossing_0_m1_write_last_time <= clock_crossing_0_m1_write;
      end if;

    end process;

    --clock_crossing_0_m1_write matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line7 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(clock_crossing_0_m1_write) /= std_logic'(clock_crossing_0_m1_write_last_time)))))) = '1' then 
          write(write_line7, now);
          write(write_line7, string'(": "));
          write(write_line7, string'("clock_crossing_0_m1_write did not heed wait!!!"));
          write(output, write_line7.all);
          deallocate (write_line7);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --clock_crossing_0_m1_writedata check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        clock_crossing_0_m1_writedata_last_time <= std_logic_vector'("00000000000000000000000000000000");
      elsif clk'event and clk = '1' then
        clock_crossing_0_m1_writedata_last_time <= clock_crossing_0_m1_writedata;
      end if;

    end process;

    --clock_crossing_0_m1_writedata matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line8 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((active_and_waiting_last_time AND to_std_logic(((clock_crossing_0_m1_writedata /= clock_crossing_0_m1_writedata_last_time)))) AND clock_crossing_0_m1_write)) = '1' then 
          write(write_line8, now);
          write(write_line8, string'(": "));
          write(write_line8, string'("clock_crossing_0_m1_writedata did not heed wait!!!"));
          write(output, write_line8.all);
          deallocate (write_line8);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity clock_crossing_0_bridge_arbitrator is 
end entity clock_crossing_0_bridge_arbitrator;


architecture europa of clock_crossing_0_bridge_arbitrator is

begin


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity rdv_fifo_for_ap_cpu_data_master_to_clock_crossing_1_s1_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC;
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity rdv_fifo_for_ap_cpu_data_master_to_clock_crossing_1_s1_module;


architecture europa of rdv_fifo_for_ap_cpu_data_master_to_clock_crossing_1_s1_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_10 :  STD_LOGIC;
                signal full_11 :  STD_LOGIC;
                signal full_12 :  STD_LOGIC;
                signal full_13 :  STD_LOGIC;
                signal full_14 :  STD_LOGIC;
                signal full_15 :  STD_LOGIC;
                signal full_16 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal full_3 :  STD_LOGIC;
                signal full_4 :  STD_LOGIC;
                signal full_5 :  STD_LOGIC;
                signal full_6 :  STD_LOGIC;
                signal full_7 :  STD_LOGIC;
                signal full_8 :  STD_LOGIC;
                signal full_9 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC;
                signal p10_full_10 :  STD_LOGIC;
                signal p10_stage_10 :  STD_LOGIC;
                signal p11_full_11 :  STD_LOGIC;
                signal p11_stage_11 :  STD_LOGIC;
                signal p12_full_12 :  STD_LOGIC;
                signal p12_stage_12 :  STD_LOGIC;
                signal p13_full_13 :  STD_LOGIC;
                signal p13_stage_13 :  STD_LOGIC;
                signal p14_full_14 :  STD_LOGIC;
                signal p14_stage_14 :  STD_LOGIC;
                signal p15_full_15 :  STD_LOGIC;
                signal p15_stage_15 :  STD_LOGIC;
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC;
                signal p2_full_2 :  STD_LOGIC;
                signal p2_stage_2 :  STD_LOGIC;
                signal p3_full_3 :  STD_LOGIC;
                signal p3_stage_3 :  STD_LOGIC;
                signal p4_full_4 :  STD_LOGIC;
                signal p4_stage_4 :  STD_LOGIC;
                signal p5_full_5 :  STD_LOGIC;
                signal p5_stage_5 :  STD_LOGIC;
                signal p6_full_6 :  STD_LOGIC;
                signal p6_stage_6 :  STD_LOGIC;
                signal p7_full_7 :  STD_LOGIC;
                signal p7_stage_7 :  STD_LOGIC;
                signal p8_full_8 :  STD_LOGIC;
                signal p8_stage_8 :  STD_LOGIC;
                signal p9_full_9 :  STD_LOGIC;
                signal p9_stage_9 :  STD_LOGIC;
                signal stage_0 :  STD_LOGIC;
                signal stage_1 :  STD_LOGIC;
                signal stage_10 :  STD_LOGIC;
                signal stage_11 :  STD_LOGIC;
                signal stage_12 :  STD_LOGIC;
                signal stage_13 :  STD_LOGIC;
                signal stage_14 :  STD_LOGIC;
                signal stage_15 :  STD_LOGIC;
                signal stage_2 :  STD_LOGIC;
                signal stage_3 :  STD_LOGIC;
                signal stage_4 :  STD_LOGIC;
                signal stage_5 :  STD_LOGIC;
                signal stage_6 :  STD_LOGIC;
                signal stage_7 :  STD_LOGIC;
                signal stage_8 :  STD_LOGIC;
                signal stage_9 :  STD_LOGIC;
                signal updated_one_count :  STD_LOGIC_VECTOR (5 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_15;
  empty <= NOT(full_0);
  full_16 <= std_logic'('0');
  --data_15, which is an e_mux
  p15_stage_15 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_16 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_15, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_15 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_15))))) = '1' then 
        if std_logic'(((sync_reset AND full_15) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_16))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_15 <= std_logic'('0');
        else
          stage_15 <= p15_stage_15;
        end if;
      end if;
    end if;

  end process;

  --control_15, which is an e_mux
  p15_full_15 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_14))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_15, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_15 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_15 <= std_logic'('0');
        else
          full_15 <= p15_full_15;
        end if;
      end if;
    end if;

  end process;

  --data_14, which is an e_mux
  p14_stage_14 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_15 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_15);
  --data_reg_14, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_14 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_14))))) = '1' then 
        if std_logic'(((sync_reset AND full_14) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_15))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_14 <= std_logic'('0');
        else
          stage_14 <= p14_stage_14;
        end if;
      end if;
    end if;

  end process;

  --control_14, which is an e_mux
  p14_full_14 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_13, full_15);
  --control_reg_14, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_14 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_14 <= std_logic'('0');
        else
          full_14 <= p14_full_14;
        end if;
      end if;
    end if;

  end process;

  --data_13, which is an e_mux
  p13_stage_13 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_14 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_14);
  --data_reg_13, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_13 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_13))))) = '1' then 
        if std_logic'(((sync_reset AND full_13) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_14))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_13 <= std_logic'('0');
        else
          stage_13 <= p13_stage_13;
        end if;
      end if;
    end if;

  end process;

  --control_13, which is an e_mux
  p13_full_13 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_12, full_14);
  --control_reg_13, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_13 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_13 <= std_logic'('0');
        else
          full_13 <= p13_full_13;
        end if;
      end if;
    end if;

  end process;

  --data_12, which is an e_mux
  p12_stage_12 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_13 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_13);
  --data_reg_12, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_12 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_12))))) = '1' then 
        if std_logic'(((sync_reset AND full_12) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_13))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_12 <= std_logic'('0');
        else
          stage_12 <= p12_stage_12;
        end if;
      end if;
    end if;

  end process;

  --control_12, which is an e_mux
  p12_full_12 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_11, full_13);
  --control_reg_12, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_12 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_12 <= std_logic'('0');
        else
          full_12 <= p12_full_12;
        end if;
      end if;
    end if;

  end process;

  --data_11, which is an e_mux
  p11_stage_11 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_12 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_12);
  --data_reg_11, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_11 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_11))))) = '1' then 
        if std_logic'(((sync_reset AND full_11) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_12))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_11 <= std_logic'('0');
        else
          stage_11 <= p11_stage_11;
        end if;
      end if;
    end if;

  end process;

  --control_11, which is an e_mux
  p11_full_11 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_10, full_12);
  --control_reg_11, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_11 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_11 <= std_logic'('0');
        else
          full_11 <= p11_full_11;
        end if;
      end if;
    end if;

  end process;

  --data_10, which is an e_mux
  p10_stage_10 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_11 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_11);
  --data_reg_10, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_10 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_10))))) = '1' then 
        if std_logic'(((sync_reset AND full_10) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_11))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_10 <= std_logic'('0');
        else
          stage_10 <= p10_stage_10;
        end if;
      end if;
    end if;

  end process;

  --control_10, which is an e_mux
  p10_full_10 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_9, full_11);
  --control_reg_10, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_10 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_10 <= std_logic'('0');
        else
          full_10 <= p10_full_10;
        end if;
      end if;
    end if;

  end process;

  --data_9, which is an e_mux
  p9_stage_9 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_10 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_10);
  --data_reg_9, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_9 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_9))))) = '1' then 
        if std_logic'(((sync_reset AND full_9) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_10))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_9 <= std_logic'('0');
        else
          stage_9 <= p9_stage_9;
        end if;
      end if;
    end if;

  end process;

  --control_9, which is an e_mux
  p9_full_9 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_8, full_10);
  --control_reg_9, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_9 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_9 <= std_logic'('0');
        else
          full_9 <= p9_full_9;
        end if;
      end if;
    end if;

  end process;

  --data_8, which is an e_mux
  p8_stage_8 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_9 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_9);
  --data_reg_8, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_8 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_8))))) = '1' then 
        if std_logic'(((sync_reset AND full_8) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_9))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_8 <= std_logic'('0');
        else
          stage_8 <= p8_stage_8;
        end if;
      end if;
    end if;

  end process;

  --control_8, which is an e_mux
  p8_full_8 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_7, full_9);
  --control_reg_8, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_8 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_8 <= std_logic'('0');
        else
          full_8 <= p8_full_8;
        end if;
      end if;
    end if;

  end process;

  --data_7, which is an e_mux
  p7_stage_7 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_8 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_8);
  --data_reg_7, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_7 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_7))))) = '1' then 
        if std_logic'(((sync_reset AND full_7) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_8))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_7 <= std_logic'('0');
        else
          stage_7 <= p7_stage_7;
        end if;
      end if;
    end if;

  end process;

  --control_7, which is an e_mux
  p7_full_7 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_6, full_8);
  --control_reg_7, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_7 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_7 <= std_logic'('0');
        else
          full_7 <= p7_full_7;
        end if;
      end if;
    end if;

  end process;

  --data_6, which is an e_mux
  p6_stage_6 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_7 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_7);
  --data_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_6 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_6))))) = '1' then 
        if std_logic'(((sync_reset AND full_6) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_7))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_6 <= std_logic'('0');
        else
          stage_6 <= p6_stage_6;
        end if;
      end if;
    end if;

  end process;

  --control_6, which is an e_mux
  p6_full_6 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_5, full_7);
  --control_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_6 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_6 <= std_logic'('0');
        else
          full_6 <= p6_full_6;
        end if;
      end if;
    end if;

  end process;

  --data_5, which is an e_mux
  p5_stage_5 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_6 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_6);
  --data_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_5))))) = '1' then 
        if std_logic'(((sync_reset AND full_5) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_6))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_5 <= std_logic'('0');
        else
          stage_5 <= p5_stage_5;
        end if;
      end if;
    end if;

  end process;

  --control_5, which is an e_mux
  p5_full_5 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_4, full_6);
  --control_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_5 <= std_logic'('0');
        else
          full_5 <= p5_full_5;
        end if;
      end if;
    end if;

  end process;

  --data_4, which is an e_mux
  p4_stage_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_5 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_5);
  --data_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_4))))) = '1' then 
        if std_logic'(((sync_reset AND full_4) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_5))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_4 <= std_logic'('0');
        else
          stage_4 <= p4_stage_4;
        end if;
      end if;
    end if;

  end process;

  --control_4, which is an e_mux
  p4_full_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_3, full_5);
  --control_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_4 <= std_logic'('0');
        else
          full_4 <= p4_full_4;
        end if;
      end if;
    end if;

  end process;

  --data_3, which is an e_mux
  p3_stage_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_4 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_4);
  --data_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_3))))) = '1' then 
        if std_logic'(((sync_reset AND full_3) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_4))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_3 <= std_logic'('0');
        else
          stage_3 <= p3_stage_3;
        end if;
      end if;
    end if;

  end process;

  --control_3, which is an e_mux
  p3_full_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_2, full_4);
  --control_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_3 <= std_logic'('0');
        else
          full_3 <= p3_full_3;
        end if;
      end if;
    end if;

  end process;

  --data_2, which is an e_mux
  p2_stage_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_3 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_3);
  --data_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_2))))) = '1' then 
        if std_logic'(((sync_reset AND full_2) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_3))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_2 <= std_logic'('0');
        else
          stage_2 <= p2_stage_2;
        end if;
      end if;
    end if;

  end process;

  --control_2, which is an e_mux
  p2_full_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_1, full_3);
  --control_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_2 <= std_logic'('0');
        else
          full_2 <= p2_full_2;
        end if;
      end if;
    end if;

  end process;

  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_2);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic'('0');
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_0, full_2);
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic'('0');
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 6);
  one_count_minus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 6);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("00000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("00000") & (A_TOSTDLOGICVECTOR(data_in))), A_WE_StdLogicVector((std_logic'(((((read AND (data_in)) AND write) AND (stage_0)))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (data_in)))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (stage_0)))) = '1'), one_count_minus_one, how_many_ones))))))), 6);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity clock_crossing_1_s1_arbitrator is 
        port (
              -- inputs:
                 signal ap_cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (25 DOWNTO 0);
                 signal ap_cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal ap_cpu_data_master_read : IN STD_LOGIC;
                 signal ap_cpu_data_master_waitrequest : IN STD_LOGIC;
                 signal ap_cpu_data_master_write : IN STD_LOGIC;
                 signal ap_cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal clk : IN STD_LOGIC;
                 signal clock_crossing_1_s1_endofpacket : IN STD_LOGIC;
                 signal clock_crossing_1_s1_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal clock_crossing_1_s1_readdatavalid : IN STD_LOGIC;
                 signal clock_crossing_1_s1_waitrequest : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal ap_cpu_data_master_granted_clock_crossing_1_s1 : OUT STD_LOGIC;
                 signal ap_cpu_data_master_qualified_request_clock_crossing_1_s1 : OUT STD_LOGIC;
                 signal ap_cpu_data_master_read_data_valid_clock_crossing_1_s1 : OUT STD_LOGIC;
                 signal ap_cpu_data_master_read_data_valid_clock_crossing_1_s1_shift_register : OUT STD_LOGIC;
                 signal ap_cpu_data_master_requests_clock_crossing_1_s1 : OUT STD_LOGIC;
                 signal clock_crossing_1_s1_address : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
                 signal clock_crossing_1_s1_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal clock_crossing_1_s1_endofpacket_from_sa : OUT STD_LOGIC;
                 signal clock_crossing_1_s1_nativeaddress : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
                 signal clock_crossing_1_s1_read : OUT STD_LOGIC;
                 signal clock_crossing_1_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal clock_crossing_1_s1_reset_n : OUT STD_LOGIC;
                 signal clock_crossing_1_s1_waitrequest_from_sa : OUT STD_LOGIC;
                 signal clock_crossing_1_s1_write : OUT STD_LOGIC;
                 signal clock_crossing_1_s1_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal d1_clock_crossing_1_s1_end_xfer : OUT STD_LOGIC
              );
end entity clock_crossing_1_s1_arbitrator;


architecture europa of clock_crossing_1_s1_arbitrator is
component rdv_fifo_for_ap_cpu_data_master_to_clock_crossing_1_s1_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC;
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component rdv_fifo_for_ap_cpu_data_master_to_clock_crossing_1_s1_module;

                signal ap_cpu_data_master_arbiterlock :  STD_LOGIC;
                signal ap_cpu_data_master_arbiterlock2 :  STD_LOGIC;
                signal ap_cpu_data_master_continuerequest :  STD_LOGIC;
                signal ap_cpu_data_master_rdv_fifo_empty_clock_crossing_1_s1 :  STD_LOGIC;
                signal ap_cpu_data_master_rdv_fifo_output_from_clock_crossing_1_s1 :  STD_LOGIC;
                signal ap_cpu_data_master_saved_grant_clock_crossing_1_s1 :  STD_LOGIC;
                signal clock_crossing_1_s1_allgrants :  STD_LOGIC;
                signal clock_crossing_1_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal clock_crossing_1_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal clock_crossing_1_s1_any_continuerequest :  STD_LOGIC;
                signal clock_crossing_1_s1_arb_counter_enable :  STD_LOGIC;
                signal clock_crossing_1_s1_arb_share_counter :  STD_LOGIC;
                signal clock_crossing_1_s1_arb_share_counter_next_value :  STD_LOGIC;
                signal clock_crossing_1_s1_arb_share_set_values :  STD_LOGIC;
                signal clock_crossing_1_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal clock_crossing_1_s1_begins_xfer :  STD_LOGIC;
                signal clock_crossing_1_s1_end_xfer :  STD_LOGIC;
                signal clock_crossing_1_s1_firsttransfer :  STD_LOGIC;
                signal clock_crossing_1_s1_grant_vector :  STD_LOGIC;
                signal clock_crossing_1_s1_in_a_read_cycle :  STD_LOGIC;
                signal clock_crossing_1_s1_in_a_write_cycle :  STD_LOGIC;
                signal clock_crossing_1_s1_master_qreq_vector :  STD_LOGIC;
                signal clock_crossing_1_s1_move_on_to_next_transaction :  STD_LOGIC;
                signal clock_crossing_1_s1_non_bursting_master_requests :  STD_LOGIC;
                signal clock_crossing_1_s1_readdatavalid_from_sa :  STD_LOGIC;
                signal clock_crossing_1_s1_reg_firsttransfer :  STD_LOGIC;
                signal clock_crossing_1_s1_slavearbiterlockenable :  STD_LOGIC;
                signal clock_crossing_1_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal clock_crossing_1_s1_unreg_firsttransfer :  STD_LOGIC;
                signal clock_crossing_1_s1_waits_for_read :  STD_LOGIC;
                signal clock_crossing_1_s1_waits_for_write :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_clock_crossing_1_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_ap_cpu_data_master_granted_clock_crossing_1_s1 :  STD_LOGIC;
                signal internal_ap_cpu_data_master_qualified_request_clock_crossing_1_s1 :  STD_LOGIC;
                signal internal_ap_cpu_data_master_read_data_valid_clock_crossing_1_s1_shift_register :  STD_LOGIC;
                signal internal_ap_cpu_data_master_requests_clock_crossing_1_s1 :  STD_LOGIC;
                signal internal_clock_crossing_1_s1_waitrequest_from_sa :  STD_LOGIC;
                signal module_input3 :  STD_LOGIC;
                signal module_input4 :  STD_LOGIC;
                signal module_input5 :  STD_LOGIC;
                signal shifted_address_to_clock_crossing_1_s1_from_ap_cpu_data_master :  STD_LOGIC_VECTOR (25 DOWNTO 0);
                signal wait_for_clock_crossing_1_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT clock_crossing_1_s1_end_xfer;
    end if;

  end process;

  clock_crossing_1_s1_begins_xfer <= NOT d1_reasons_to_wait AND (internal_ap_cpu_data_master_qualified_request_clock_crossing_1_s1);
  --assign clock_crossing_1_s1_readdata_from_sa = clock_crossing_1_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  clock_crossing_1_s1_readdata_from_sa <= clock_crossing_1_s1_readdata;
  internal_ap_cpu_data_master_requests_clock_crossing_1_s1 <= to_std_logic(((Std_Logic_Vector'(ap_cpu_data_master_address_to_slave(25 DOWNTO 8) & std_logic_vector'("00000000")) = std_logic_vector'("01000000000000000000000000")))) AND ((ap_cpu_data_master_read OR ap_cpu_data_master_write));
  --assign clock_crossing_1_s1_waitrequest_from_sa = clock_crossing_1_s1_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_clock_crossing_1_s1_waitrequest_from_sa <= clock_crossing_1_s1_waitrequest;
  --assign clock_crossing_1_s1_readdatavalid_from_sa = clock_crossing_1_s1_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  clock_crossing_1_s1_readdatavalid_from_sa <= clock_crossing_1_s1_readdatavalid;
  --clock_crossing_1_s1_arb_share_counter set values, which is an e_mux
  clock_crossing_1_s1_arb_share_set_values <= std_logic'('1');
  --clock_crossing_1_s1_non_bursting_master_requests mux, which is an e_mux
  clock_crossing_1_s1_non_bursting_master_requests <= internal_ap_cpu_data_master_requests_clock_crossing_1_s1;
  --clock_crossing_1_s1_any_bursting_master_saved_grant mux, which is an e_mux
  clock_crossing_1_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --clock_crossing_1_s1_arb_share_counter_next_value assignment, which is an e_assign
  clock_crossing_1_s1_arb_share_counter_next_value <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(clock_crossing_1_s1_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(clock_crossing_1_s1_arb_share_set_values))) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(clock_crossing_1_s1_arb_share_counter) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(clock_crossing_1_s1_arb_share_counter))) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))));
  --clock_crossing_1_s1_allgrants all slave grants, which is an e_mux
  clock_crossing_1_s1_allgrants <= clock_crossing_1_s1_grant_vector;
  --clock_crossing_1_s1_end_xfer assignment, which is an e_assign
  clock_crossing_1_s1_end_xfer <= NOT ((clock_crossing_1_s1_waits_for_read OR clock_crossing_1_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_clock_crossing_1_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_clock_crossing_1_s1 <= clock_crossing_1_s1_end_xfer AND (((NOT clock_crossing_1_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --clock_crossing_1_s1_arb_share_counter arbitration counter enable, which is an e_assign
  clock_crossing_1_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_clock_crossing_1_s1 AND clock_crossing_1_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_clock_crossing_1_s1 AND NOT clock_crossing_1_s1_non_bursting_master_requests));
  --clock_crossing_1_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      clock_crossing_1_s1_arb_share_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(clock_crossing_1_s1_arb_counter_enable) = '1' then 
        clock_crossing_1_s1_arb_share_counter <= clock_crossing_1_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --clock_crossing_1_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      clock_crossing_1_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clock_crossing_1_s1_master_qreq_vector AND end_xfer_arb_share_counter_term_clock_crossing_1_s1)) OR ((end_xfer_arb_share_counter_term_clock_crossing_1_s1 AND NOT clock_crossing_1_s1_non_bursting_master_requests)))) = '1' then 
        clock_crossing_1_s1_slavearbiterlockenable <= clock_crossing_1_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --ap_cpu/data_master clock_crossing_1/s1 arbiterlock, which is an e_assign
  ap_cpu_data_master_arbiterlock <= clock_crossing_1_s1_slavearbiterlockenable AND ap_cpu_data_master_continuerequest;
  --clock_crossing_1_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  clock_crossing_1_s1_slavearbiterlockenable2 <= clock_crossing_1_s1_arb_share_counter_next_value;
  --ap_cpu/data_master clock_crossing_1/s1 arbiterlock2, which is an e_assign
  ap_cpu_data_master_arbiterlock2 <= clock_crossing_1_s1_slavearbiterlockenable2 AND ap_cpu_data_master_continuerequest;
  --clock_crossing_1_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  clock_crossing_1_s1_any_continuerequest <= std_logic'('1');
  --ap_cpu_data_master_continuerequest continued request, which is an e_assign
  ap_cpu_data_master_continuerequest <= std_logic'('1');
  internal_ap_cpu_data_master_qualified_request_clock_crossing_1_s1 <= internal_ap_cpu_data_master_requests_clock_crossing_1_s1 AND NOT ((((ap_cpu_data_master_read AND ((NOT ap_cpu_data_master_waitrequest OR (internal_ap_cpu_data_master_read_data_valid_clock_crossing_1_s1_shift_register))))) OR (((NOT ap_cpu_data_master_waitrequest) AND ap_cpu_data_master_write))));
  --unique name for clock_crossing_1_s1_move_on_to_next_transaction, which is an e_assign
  clock_crossing_1_s1_move_on_to_next_transaction <= clock_crossing_1_s1_readdatavalid_from_sa;
  --rdv_fifo_for_ap_cpu_data_master_to_clock_crossing_1_s1, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_ap_cpu_data_master_to_clock_crossing_1_s1 : rdv_fifo_for_ap_cpu_data_master_to_clock_crossing_1_s1_module
    port map(
      data_out => ap_cpu_data_master_rdv_fifo_output_from_clock_crossing_1_s1,
      empty => open,
      fifo_contains_ones_n => ap_cpu_data_master_rdv_fifo_empty_clock_crossing_1_s1,
      full => open,
      clear_fifo => module_input3,
      clk => clk,
      data_in => internal_ap_cpu_data_master_granted_clock_crossing_1_s1,
      read => clock_crossing_1_s1_move_on_to_next_transaction,
      reset_n => reset_n,
      sync_reset => module_input4,
      write => module_input5
    );

  module_input3 <= std_logic'('0');
  module_input4 <= std_logic'('0');
  module_input5 <= in_a_read_cycle AND NOT clock_crossing_1_s1_waits_for_read;

  internal_ap_cpu_data_master_read_data_valid_clock_crossing_1_s1_shift_register <= NOT ap_cpu_data_master_rdv_fifo_empty_clock_crossing_1_s1;
  --local readdatavalid ap_cpu_data_master_read_data_valid_clock_crossing_1_s1, which is an e_mux
  ap_cpu_data_master_read_data_valid_clock_crossing_1_s1 <= clock_crossing_1_s1_readdatavalid_from_sa;
  --clock_crossing_1_s1_writedata mux, which is an e_mux
  clock_crossing_1_s1_writedata <= ap_cpu_data_master_writedata;
  --assign clock_crossing_1_s1_endofpacket_from_sa = clock_crossing_1_s1_endofpacket so that symbol knows where to group signals which may go to master only, which is an e_assign
  clock_crossing_1_s1_endofpacket_from_sa <= clock_crossing_1_s1_endofpacket;
  --master is always granted when requested
  internal_ap_cpu_data_master_granted_clock_crossing_1_s1 <= internal_ap_cpu_data_master_qualified_request_clock_crossing_1_s1;
  --ap_cpu/data_master saved-grant clock_crossing_1/s1, which is an e_assign
  ap_cpu_data_master_saved_grant_clock_crossing_1_s1 <= internal_ap_cpu_data_master_requests_clock_crossing_1_s1;
  --allow new arb cycle for clock_crossing_1/s1, which is an e_assign
  clock_crossing_1_s1_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  clock_crossing_1_s1_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  clock_crossing_1_s1_master_qreq_vector <= std_logic'('1');
  --clock_crossing_1_s1_reset_n assignment, which is an e_assign
  clock_crossing_1_s1_reset_n <= reset_n;
  --clock_crossing_1_s1_firsttransfer first transaction, which is an e_assign
  clock_crossing_1_s1_firsttransfer <= A_WE_StdLogic((std_logic'(clock_crossing_1_s1_begins_xfer) = '1'), clock_crossing_1_s1_unreg_firsttransfer, clock_crossing_1_s1_reg_firsttransfer);
  --clock_crossing_1_s1_unreg_firsttransfer first transaction, which is an e_assign
  clock_crossing_1_s1_unreg_firsttransfer <= NOT ((clock_crossing_1_s1_slavearbiterlockenable AND clock_crossing_1_s1_any_continuerequest));
  --clock_crossing_1_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      clock_crossing_1_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(clock_crossing_1_s1_begins_xfer) = '1' then 
        clock_crossing_1_s1_reg_firsttransfer <= clock_crossing_1_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --clock_crossing_1_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  clock_crossing_1_s1_beginbursttransfer_internal <= clock_crossing_1_s1_begins_xfer;
  --clock_crossing_1_s1_read assignment, which is an e_mux
  clock_crossing_1_s1_read <= internal_ap_cpu_data_master_granted_clock_crossing_1_s1 AND ap_cpu_data_master_read;
  --clock_crossing_1_s1_write assignment, which is an e_mux
  clock_crossing_1_s1_write <= internal_ap_cpu_data_master_granted_clock_crossing_1_s1 AND ap_cpu_data_master_write;
  shifted_address_to_clock_crossing_1_s1_from_ap_cpu_data_master <= ap_cpu_data_master_address_to_slave;
  --clock_crossing_1_s1_address mux, which is an e_mux
  clock_crossing_1_s1_address <= A_EXT (A_SRL(shifted_address_to_clock_crossing_1_s1_from_ap_cpu_data_master,std_logic_vector'("00000000000000000000000000000010")), 6);
  --slaveid clock_crossing_1_s1_nativeaddress nativeaddress mux, which is an e_mux
  clock_crossing_1_s1_nativeaddress <= A_EXT (A_SRL(ap_cpu_data_master_address_to_slave,std_logic_vector'("00000000000000000000000000000010")), 6);
  --d1_clock_crossing_1_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_clock_crossing_1_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_clock_crossing_1_s1_end_xfer <= clock_crossing_1_s1_end_xfer;
    end if;

  end process;

  --clock_crossing_1_s1_waits_for_read in a cycle, which is an e_mux
  clock_crossing_1_s1_waits_for_read <= clock_crossing_1_s1_in_a_read_cycle AND internal_clock_crossing_1_s1_waitrequest_from_sa;
  --clock_crossing_1_s1_in_a_read_cycle assignment, which is an e_assign
  clock_crossing_1_s1_in_a_read_cycle <= internal_ap_cpu_data_master_granted_clock_crossing_1_s1 AND ap_cpu_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= clock_crossing_1_s1_in_a_read_cycle;
  --clock_crossing_1_s1_waits_for_write in a cycle, which is an e_mux
  clock_crossing_1_s1_waits_for_write <= clock_crossing_1_s1_in_a_write_cycle AND internal_clock_crossing_1_s1_waitrequest_from_sa;
  --clock_crossing_1_s1_in_a_write_cycle assignment, which is an e_assign
  clock_crossing_1_s1_in_a_write_cycle <= internal_ap_cpu_data_master_granted_clock_crossing_1_s1 AND ap_cpu_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= clock_crossing_1_s1_in_a_write_cycle;
  wait_for_clock_crossing_1_s1_counter <= std_logic'('0');
  --clock_crossing_1_s1_byteenable byte enable port mux, which is an e_mux
  clock_crossing_1_s1_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_ap_cpu_data_master_granted_clock_crossing_1_s1)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (ap_cpu_data_master_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))), 4);
  --vhdl renameroo for output signals
  ap_cpu_data_master_granted_clock_crossing_1_s1 <= internal_ap_cpu_data_master_granted_clock_crossing_1_s1;
  --vhdl renameroo for output signals
  ap_cpu_data_master_qualified_request_clock_crossing_1_s1 <= internal_ap_cpu_data_master_qualified_request_clock_crossing_1_s1;
  --vhdl renameroo for output signals
  ap_cpu_data_master_read_data_valid_clock_crossing_1_s1_shift_register <= internal_ap_cpu_data_master_read_data_valid_clock_crossing_1_s1_shift_register;
  --vhdl renameroo for output signals
  ap_cpu_data_master_requests_clock_crossing_1_s1 <= internal_ap_cpu_data_master_requests_clock_crossing_1_s1;
  --vhdl renameroo for output signals
  clock_crossing_1_s1_waitrequest_from_sa <= internal_clock_crossing_1_s1_waitrequest_from_sa;
--synthesis translate_off
    --clock_crossing_1/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity clock_crossing_1_m1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal clock_crossing_1_m1_address : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal clock_crossing_1_m1_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal clock_crossing_1_m1_granted_digio_pio_s1 : IN STD_LOGIC;
                 signal clock_crossing_1_m1_granted_node_switch_pio_s1 : IN STD_LOGIC;
                 signal clock_crossing_1_m1_granted_portconf_pio_s1 : IN STD_LOGIC;
                 signal clock_crossing_1_m1_granted_sync_irq_s1 : IN STD_LOGIC;
                 signal clock_crossing_1_m1_granted_sysid_control_slave : IN STD_LOGIC;
                 signal clock_crossing_1_m1_granted_system_timer_ap_s1 : IN STD_LOGIC;
                 signal clock_crossing_1_m1_qualified_request_digio_pio_s1 : IN STD_LOGIC;
                 signal clock_crossing_1_m1_qualified_request_node_switch_pio_s1 : IN STD_LOGIC;
                 signal clock_crossing_1_m1_qualified_request_portconf_pio_s1 : IN STD_LOGIC;
                 signal clock_crossing_1_m1_qualified_request_sync_irq_s1 : IN STD_LOGIC;
                 signal clock_crossing_1_m1_qualified_request_sysid_control_slave : IN STD_LOGIC;
                 signal clock_crossing_1_m1_qualified_request_system_timer_ap_s1 : IN STD_LOGIC;
                 signal clock_crossing_1_m1_read : IN STD_LOGIC;
                 signal clock_crossing_1_m1_read_data_valid_digio_pio_s1 : IN STD_LOGIC;
                 signal clock_crossing_1_m1_read_data_valid_node_switch_pio_s1 : IN STD_LOGIC;
                 signal clock_crossing_1_m1_read_data_valid_portconf_pio_s1 : IN STD_LOGIC;
                 signal clock_crossing_1_m1_read_data_valid_sync_irq_s1 : IN STD_LOGIC;
                 signal clock_crossing_1_m1_read_data_valid_sysid_control_slave : IN STD_LOGIC;
                 signal clock_crossing_1_m1_read_data_valid_system_timer_ap_s1 : IN STD_LOGIC;
                 signal clock_crossing_1_m1_requests_digio_pio_s1 : IN STD_LOGIC;
                 signal clock_crossing_1_m1_requests_node_switch_pio_s1 : IN STD_LOGIC;
                 signal clock_crossing_1_m1_requests_portconf_pio_s1 : IN STD_LOGIC;
                 signal clock_crossing_1_m1_requests_sync_irq_s1 : IN STD_LOGIC;
                 signal clock_crossing_1_m1_requests_sysid_control_slave : IN STD_LOGIC;
                 signal clock_crossing_1_m1_requests_system_timer_ap_s1 : IN STD_LOGIC;
                 signal clock_crossing_1_m1_write : IN STD_LOGIC;
                 signal clock_crossing_1_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal d1_digio_pio_s1_end_xfer : IN STD_LOGIC;
                 signal d1_node_switch_pio_s1_end_xfer : IN STD_LOGIC;
                 signal d1_portconf_pio_s1_end_xfer : IN STD_LOGIC;
                 signal d1_sync_irq_s1_end_xfer : IN STD_LOGIC;
                 signal d1_sysid_control_slave_end_xfer : IN STD_LOGIC;
                 signal d1_system_timer_ap_s1_end_xfer : IN STD_LOGIC;
                 signal digio_pio_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal node_switch_pio_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal portconf_pio_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;
                 signal sync_irq_s1_readdata_from_sa : IN STD_LOGIC;
                 signal sysid_control_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal system_timer_ap_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

              -- outputs:
                 signal clock_crossing_1_m1_address_to_slave : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal clock_crossing_1_m1_latency_counter : OUT STD_LOGIC;
                 signal clock_crossing_1_m1_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal clock_crossing_1_m1_readdatavalid : OUT STD_LOGIC;
                 signal clock_crossing_1_m1_reset_n : OUT STD_LOGIC;
                 signal clock_crossing_1_m1_waitrequest : OUT STD_LOGIC
              );
end entity clock_crossing_1_m1_arbitrator;


architecture europa of clock_crossing_1_m1_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal clock_crossing_1_m1_address_last_time :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal clock_crossing_1_m1_byteenable_last_time :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal clock_crossing_1_m1_is_granted_some_slave :  STD_LOGIC;
                signal clock_crossing_1_m1_read_but_no_slave_selected :  STD_LOGIC;
                signal clock_crossing_1_m1_read_last_time :  STD_LOGIC;
                signal clock_crossing_1_m1_run :  STD_LOGIC;
                signal clock_crossing_1_m1_write_last_time :  STD_LOGIC;
                signal clock_crossing_1_m1_writedata_last_time :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal internal_clock_crossing_1_m1_address_to_slave :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal internal_clock_crossing_1_m1_latency_counter :  STD_LOGIC;
                signal internal_clock_crossing_1_m1_waitrequest :  STD_LOGIC;
                signal latency_load_value :  STD_LOGIC;
                signal p1_clock_crossing_1_m1_latency_counter :  STD_LOGIC;
                signal pre_flush_clock_crossing_1_m1_readdatavalid :  STD_LOGIC;
                signal r_0 :  STD_LOGIC;
                signal r_1 :  STD_LOGIC;
                signal r_2 :  STD_LOGIC;

begin

  --r_0 master_run cascaded wait assignment, which is an e_assign
  r_0 <= Vector_To_Std_Logic((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((clock_crossing_1_m1_qualified_request_digio_pio_s1 OR NOT clock_crossing_1_m1_requests_digio_pio_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT clock_crossing_1_m1_qualified_request_digio_pio_s1 OR NOT clock_crossing_1_m1_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT d1_digio_pio_s1_end_xfer)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(clock_crossing_1_m1_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT clock_crossing_1_m1_qualified_request_digio_pio_s1 OR NOT clock_crossing_1_m1_write)))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(clock_crossing_1_m1_write)))))))));
  --cascaded wait assignment, which is an e_assign
  clock_crossing_1_m1_run <= (r_0 AND r_1) AND r_2;
  --r_1 master_run cascaded wait assignment, which is an e_assign
  r_1 <= Vector_To_Std_Logic((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((clock_crossing_1_m1_qualified_request_node_switch_pio_s1 OR NOT clock_crossing_1_m1_requests_node_switch_pio_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT clock_crossing_1_m1_qualified_request_node_switch_pio_s1 OR NOT clock_crossing_1_m1_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT d1_node_switch_pio_s1_end_xfer)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(clock_crossing_1_m1_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT clock_crossing_1_m1_qualified_request_node_switch_pio_s1 OR NOT clock_crossing_1_m1_write)))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(clock_crossing_1_m1_write)))))))));
  --r_2 master_run cascaded wait assignment, which is an e_assign
  r_2 <= Vector_To_Std_Logic(((((((((((((((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((clock_crossing_1_m1_qualified_request_portconf_pio_s1 OR NOT clock_crossing_1_m1_requests_portconf_pio_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT clock_crossing_1_m1_qualified_request_portconf_pio_s1 OR NOT clock_crossing_1_m1_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT d1_portconf_pio_s1_end_xfer)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(clock_crossing_1_m1_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT clock_crossing_1_m1_qualified_request_portconf_pio_s1 OR NOT clock_crossing_1_m1_write)))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(clock_crossing_1_m1_write)))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((clock_crossing_1_m1_qualified_request_sync_irq_s1 OR NOT clock_crossing_1_m1_requests_sync_irq_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT clock_crossing_1_m1_qualified_request_sync_irq_s1 OR NOT clock_crossing_1_m1_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT d1_sync_irq_s1_end_xfer)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(clock_crossing_1_m1_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT clock_crossing_1_m1_qualified_request_sync_irq_s1 OR NOT clock_crossing_1_m1_write)))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(clock_crossing_1_m1_write)))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((clock_crossing_1_m1_qualified_request_sysid_control_slave OR NOT clock_crossing_1_m1_requests_sysid_control_slave)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((clock_crossing_1_m1_granted_sysid_control_slave OR NOT clock_crossing_1_m1_qualified_request_sysid_control_slave)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT clock_crossing_1_m1_qualified_request_sysid_control_slave OR NOT clock_crossing_1_m1_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT d1_sysid_control_slave_end_xfer)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(clock_crossing_1_m1_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT clock_crossing_1_m1_qualified_request_sysid_control_slave OR NOT clock_crossing_1_m1_write)))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(clock_crossing_1_m1_write)))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((clock_crossing_1_m1_qualified_request_system_timer_ap_s1 OR NOT clock_crossing_1_m1_requests_system_timer_ap_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT clock_crossing_1_m1_qualified_request_system_timer_ap_s1 OR NOT clock_crossing_1_m1_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT d1_system_timer_ap_s1_end_xfer)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(clock_crossing_1_m1_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT clock_crossing_1_m1_qualified_request_system_timer_ap_s1 OR NOT clock_crossing_1_m1_write)))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(clock_crossing_1_m1_write)))))))));
  --optimize select-logic by passing only those address bits which matter.
  internal_clock_crossing_1_m1_address_to_slave <= clock_crossing_1_m1_address(7 DOWNTO 0);
  --clock_crossing_1_m1_read_but_no_slave_selected assignment, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      clock_crossing_1_m1_read_but_no_slave_selected <= std_logic'('0');
    elsif clk'event and clk = '1' then
      clock_crossing_1_m1_read_but_no_slave_selected <= (clock_crossing_1_m1_read AND clock_crossing_1_m1_run) AND NOT clock_crossing_1_m1_is_granted_some_slave;
    end if;

  end process;

  --some slave is getting selected, which is an e_mux
  clock_crossing_1_m1_is_granted_some_slave <= ((((clock_crossing_1_m1_granted_digio_pio_s1 OR clock_crossing_1_m1_granted_node_switch_pio_s1) OR clock_crossing_1_m1_granted_portconf_pio_s1) OR clock_crossing_1_m1_granted_sync_irq_s1) OR clock_crossing_1_m1_granted_sysid_control_slave) OR clock_crossing_1_m1_granted_system_timer_ap_s1;
  --latent slave read data valids which may be flushed, which is an e_mux
  pre_flush_clock_crossing_1_m1_readdatavalid <= std_logic'('0');
  --latent slave read data valid which is not flushed, which is an e_mux
  clock_crossing_1_m1_readdatavalid <= ((((((((((((((((clock_crossing_1_m1_read_but_no_slave_selected OR pre_flush_clock_crossing_1_m1_readdatavalid) OR clock_crossing_1_m1_read_data_valid_digio_pio_s1) OR clock_crossing_1_m1_read_but_no_slave_selected) OR pre_flush_clock_crossing_1_m1_readdatavalid) OR clock_crossing_1_m1_read_data_valid_node_switch_pio_s1) OR clock_crossing_1_m1_read_but_no_slave_selected) OR pre_flush_clock_crossing_1_m1_readdatavalid) OR clock_crossing_1_m1_read_data_valid_portconf_pio_s1) OR clock_crossing_1_m1_read_but_no_slave_selected) OR pre_flush_clock_crossing_1_m1_readdatavalid) OR clock_crossing_1_m1_read_data_valid_sync_irq_s1) OR clock_crossing_1_m1_read_but_no_slave_selected) OR pre_flush_clock_crossing_1_m1_readdatavalid) OR clock_crossing_1_m1_read_data_valid_sysid_control_slave) OR clock_crossing_1_m1_read_but_no_slave_selected) OR pre_flush_clock_crossing_1_m1_readdatavalid) OR clock_crossing_1_m1_read_data_valid_system_timer_ap_s1;
  --clock_crossing_1/m1 readdata mux, which is an e_mux
  clock_crossing_1_m1_readdata <= ((((((A_REP(NOT ((clock_crossing_1_m1_qualified_request_digio_pio_s1 AND clock_crossing_1_m1_read)) , 32) OR digio_pio_s1_readdata_from_sa)) AND ((A_REP(NOT ((clock_crossing_1_m1_qualified_request_node_switch_pio_s1 AND clock_crossing_1_m1_read)) , 32) OR (std_logic_vector'("000000000000000000000000") & (node_switch_pio_s1_readdata_from_sa))))) AND ((A_REP(NOT ((clock_crossing_1_m1_qualified_request_portconf_pio_s1 AND clock_crossing_1_m1_read)) , 32) OR (std_logic_vector'("0000000000000000000000000000") & (portconf_pio_s1_readdata_from_sa))))) AND ((A_REP(NOT ((clock_crossing_1_m1_qualified_request_sync_irq_s1 AND clock_crossing_1_m1_read)) , 32) OR (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(sync_irq_s1_readdata_from_sa)))))) AND ((A_REP(NOT ((clock_crossing_1_m1_qualified_request_sysid_control_slave AND clock_crossing_1_m1_read)) , 32) OR sysid_control_slave_readdata_from_sa))) AND ((A_REP(NOT ((clock_crossing_1_m1_qualified_request_system_timer_ap_s1 AND clock_crossing_1_m1_read)) , 32) OR (std_logic_vector'("0000000000000000") & (system_timer_ap_s1_readdata_from_sa))));
  --actual waitrequest port, which is an e_assign
  internal_clock_crossing_1_m1_waitrequest <= NOT clock_crossing_1_m1_run;
  --latent max counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      internal_clock_crossing_1_m1_latency_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      internal_clock_crossing_1_m1_latency_counter <= p1_clock_crossing_1_m1_latency_counter;
    end if;

  end process;

  --latency counter load mux, which is an e_mux
  p1_clock_crossing_1_m1_latency_counter <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(((clock_crossing_1_m1_run AND clock_crossing_1_m1_read))) = '1'), (std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(latency_load_value))), A_WE_StdLogicVector((std_logic'((internal_clock_crossing_1_m1_latency_counter)) = '1'), ((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(internal_clock_crossing_1_m1_latency_counter))) - std_logic_vector'("000000000000000000000000000000001")), std_logic_vector'("000000000000000000000000000000000"))));
  --read latency load values, which is an e_mux
  latency_load_value <= std_logic'('0');
  --clock_crossing_1_m1_reset_n assignment, which is an e_assign
  clock_crossing_1_m1_reset_n <= reset_n;
  --vhdl renameroo for output signals
  clock_crossing_1_m1_address_to_slave <= internal_clock_crossing_1_m1_address_to_slave;
  --vhdl renameroo for output signals
  clock_crossing_1_m1_latency_counter <= internal_clock_crossing_1_m1_latency_counter;
  --vhdl renameroo for output signals
  clock_crossing_1_m1_waitrequest <= internal_clock_crossing_1_m1_waitrequest;
--synthesis translate_off
    --clock_crossing_1_m1_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        clock_crossing_1_m1_address_last_time <= std_logic_vector'("00000000");
      elsif clk'event and clk = '1' then
        clock_crossing_1_m1_address_last_time <= clock_crossing_1_m1_address;
      end if;

    end process;

    --clock_crossing_1/m1 waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_clock_crossing_1_m1_waitrequest AND ((clock_crossing_1_m1_read OR clock_crossing_1_m1_write));
      end if;

    end process;

    --clock_crossing_1_m1_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line9 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((clock_crossing_1_m1_address /= clock_crossing_1_m1_address_last_time))))) = '1' then 
          write(write_line9, now);
          write(write_line9, string'(": "));
          write(write_line9, string'("clock_crossing_1_m1_address did not heed wait!!!"));
          write(output, write_line9.all);
          deallocate (write_line9);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --clock_crossing_1_m1_byteenable check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        clock_crossing_1_m1_byteenable_last_time <= std_logic_vector'("0000");
      elsif clk'event and clk = '1' then
        clock_crossing_1_m1_byteenable_last_time <= clock_crossing_1_m1_byteenable;
      end if;

    end process;

    --clock_crossing_1_m1_byteenable matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line10 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((clock_crossing_1_m1_byteenable /= clock_crossing_1_m1_byteenable_last_time))))) = '1' then 
          write(write_line10, now);
          write(write_line10, string'(": "));
          write(write_line10, string'("clock_crossing_1_m1_byteenable did not heed wait!!!"));
          write(output, write_line10.all);
          deallocate (write_line10);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --clock_crossing_1_m1_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        clock_crossing_1_m1_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        clock_crossing_1_m1_read_last_time <= clock_crossing_1_m1_read;
      end if;

    end process;

    --clock_crossing_1_m1_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line11 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(clock_crossing_1_m1_read) /= std_logic'(clock_crossing_1_m1_read_last_time)))))) = '1' then 
          write(write_line11, now);
          write(write_line11, string'(": "));
          write(write_line11, string'("clock_crossing_1_m1_read did not heed wait!!!"));
          write(output, write_line11.all);
          deallocate (write_line11);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --clock_crossing_1_m1_write check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        clock_crossing_1_m1_write_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        clock_crossing_1_m1_write_last_time <= clock_crossing_1_m1_write;
      end if;

    end process;

    --clock_crossing_1_m1_write matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line12 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(clock_crossing_1_m1_write) /= std_logic'(clock_crossing_1_m1_write_last_time)))))) = '1' then 
          write(write_line12, now);
          write(write_line12, string'(": "));
          write(write_line12, string'("clock_crossing_1_m1_write did not heed wait!!!"));
          write(output, write_line12.all);
          deallocate (write_line12);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --clock_crossing_1_m1_writedata check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        clock_crossing_1_m1_writedata_last_time <= std_logic_vector'("00000000000000000000000000000000");
      elsif clk'event and clk = '1' then
        clock_crossing_1_m1_writedata_last_time <= clock_crossing_1_m1_writedata;
      end if;

    end process;

    --clock_crossing_1_m1_writedata matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line13 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((active_and_waiting_last_time AND to_std_logic(((clock_crossing_1_m1_writedata /= clock_crossing_1_m1_writedata_last_time)))) AND clock_crossing_1_m1_write)) = '1' then 
          write(write_line13, now);
          write(write_line13, string'(": "));
          write(write_line13, string'("clock_crossing_1_m1_writedata did not heed wait!!!"));
          write(output, write_line13.all);
          deallocate (write_line13);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity clock_crossing_1_bridge_arbitrator is 
end entity clock_crossing_1_bridge_arbitrator;


architecture europa of clock_crossing_1_bridge_arbitrator is

begin


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity cnApi_Av2Av_0_ap_arbitrator is 
        port (
              -- inputs:
                 signal ap_cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (25 DOWNTO 0);
                 signal ap_cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal ap_cpu_data_master_read : IN STD_LOGIC;
                 signal ap_cpu_data_master_waitrequest : IN STD_LOGIC;
                 signal ap_cpu_data_master_write : IN STD_LOGIC;
                 signal ap_cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal clk : IN STD_LOGIC;
                 signal cnApi_Av2Av_0_ap_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal ap_cpu_data_master_granted_cnApi_Av2Av_0_ap : OUT STD_LOGIC;
                 signal ap_cpu_data_master_qualified_request_cnApi_Av2Av_0_ap : OUT STD_LOGIC;
                 signal ap_cpu_data_master_read_data_valid_cnApi_Av2Av_0_ap : OUT STD_LOGIC;
                 signal ap_cpu_data_master_requests_cnApi_Av2Av_0_ap : OUT STD_LOGIC;
                 signal cnApi_Av2Av_0_ap_address : OUT STD_LOGIC_VECTOR (14 DOWNTO 0);
                 signal cnApi_Av2Av_0_ap_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cnApi_Av2Av_0_ap_chipselect : OUT STD_LOGIC;
                 signal cnApi_Av2Av_0_ap_read : OUT STD_LOGIC;
                 signal cnApi_Av2Av_0_ap_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal cnApi_Av2Av_0_ap_reset : OUT STD_LOGIC;
                 signal cnApi_Av2Av_0_ap_wait_counter_eq_0 : OUT STD_LOGIC;
                 signal cnApi_Av2Av_0_ap_write : OUT STD_LOGIC;
                 signal cnApi_Av2Av_0_ap_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal d1_cnApi_Av2Av_0_ap_end_xfer : OUT STD_LOGIC
              );
end entity cnApi_Av2Av_0_ap_arbitrator;


architecture europa of cnApi_Av2Av_0_ap_arbitrator is
                signal ap_cpu_data_master_arbiterlock :  STD_LOGIC;
                signal ap_cpu_data_master_arbiterlock2 :  STD_LOGIC;
                signal ap_cpu_data_master_continuerequest :  STD_LOGIC;
                signal ap_cpu_data_master_saved_grant_cnApi_Av2Av_0_ap :  STD_LOGIC;
                signal cnApi_Av2Av_0_ap_allgrants :  STD_LOGIC;
                signal cnApi_Av2Av_0_ap_allow_new_arb_cycle :  STD_LOGIC;
                signal cnApi_Av2Av_0_ap_any_bursting_master_saved_grant :  STD_LOGIC;
                signal cnApi_Av2Av_0_ap_any_continuerequest :  STD_LOGIC;
                signal cnApi_Av2Av_0_ap_arb_counter_enable :  STD_LOGIC;
                signal cnApi_Av2Av_0_ap_arb_share_counter :  STD_LOGIC;
                signal cnApi_Av2Av_0_ap_arb_share_counter_next_value :  STD_LOGIC;
                signal cnApi_Av2Av_0_ap_arb_share_set_values :  STD_LOGIC;
                signal cnApi_Av2Av_0_ap_beginbursttransfer_internal :  STD_LOGIC;
                signal cnApi_Av2Av_0_ap_begins_xfer :  STD_LOGIC;
                signal cnApi_Av2Av_0_ap_counter_load_value :  STD_LOGIC;
                signal cnApi_Av2Av_0_ap_end_xfer :  STD_LOGIC;
                signal cnApi_Av2Av_0_ap_firsttransfer :  STD_LOGIC;
                signal cnApi_Av2Av_0_ap_grant_vector :  STD_LOGIC;
                signal cnApi_Av2Av_0_ap_in_a_read_cycle :  STD_LOGIC;
                signal cnApi_Av2Av_0_ap_in_a_write_cycle :  STD_LOGIC;
                signal cnApi_Av2Av_0_ap_master_qreq_vector :  STD_LOGIC;
                signal cnApi_Av2Av_0_ap_non_bursting_master_requests :  STD_LOGIC;
                signal cnApi_Av2Av_0_ap_reg_firsttransfer :  STD_LOGIC;
                signal cnApi_Av2Av_0_ap_slavearbiterlockenable :  STD_LOGIC;
                signal cnApi_Av2Av_0_ap_slavearbiterlockenable2 :  STD_LOGIC;
                signal cnApi_Av2Av_0_ap_unreg_firsttransfer :  STD_LOGIC;
                signal cnApi_Av2Av_0_ap_wait_counter :  STD_LOGIC;
                signal cnApi_Av2Av_0_ap_waits_for_read :  STD_LOGIC;
                signal cnApi_Av2Av_0_ap_waits_for_write :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_cnApi_Av2Av_0_ap :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_ap_cpu_data_master_granted_cnApi_Av2Av_0_ap :  STD_LOGIC;
                signal internal_ap_cpu_data_master_qualified_request_cnApi_Av2Av_0_ap :  STD_LOGIC;
                signal internal_ap_cpu_data_master_requests_cnApi_Av2Av_0_ap :  STD_LOGIC;
                signal internal_cnApi_Av2Av_0_ap_wait_counter_eq_0 :  STD_LOGIC;
                signal shifted_address_to_cnApi_Av2Av_0_ap_from_ap_cpu_data_master :  STD_LOGIC_VECTOR (25 DOWNTO 0);
                signal wait_for_cnApi_Av2Av_0_ap_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT cnApi_Av2Av_0_ap_end_xfer;
    end if;

  end process;

  cnApi_Av2Av_0_ap_begins_xfer <= NOT d1_reasons_to_wait AND (internal_ap_cpu_data_master_qualified_request_cnApi_Av2Av_0_ap);
  --assign cnApi_Av2Av_0_ap_readdata_from_sa = cnApi_Av2Av_0_ap_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  cnApi_Av2Av_0_ap_readdata_from_sa <= cnApi_Av2Av_0_ap_readdata;
  internal_ap_cpu_data_master_requests_cnApi_Av2Av_0_ap <= to_std_logic(((Std_Logic_Vector'(ap_cpu_data_master_address_to_slave(25 DOWNTO 17) & std_logic_vector'("00000000000000000")) = std_logic_vector'("11000000000000000000000000")))) AND ((ap_cpu_data_master_read OR ap_cpu_data_master_write));
  --cnApi_Av2Av_0_ap_arb_share_counter set values, which is an e_mux
  cnApi_Av2Av_0_ap_arb_share_set_values <= std_logic'('1');
  --cnApi_Av2Av_0_ap_non_bursting_master_requests mux, which is an e_mux
  cnApi_Av2Av_0_ap_non_bursting_master_requests <= internal_ap_cpu_data_master_requests_cnApi_Av2Av_0_ap;
  --cnApi_Av2Av_0_ap_any_bursting_master_saved_grant mux, which is an e_mux
  cnApi_Av2Av_0_ap_any_bursting_master_saved_grant <= std_logic'('0');
  --cnApi_Av2Av_0_ap_arb_share_counter_next_value assignment, which is an e_assign
  cnApi_Av2Av_0_ap_arb_share_counter_next_value <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(cnApi_Av2Av_0_ap_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cnApi_Av2Av_0_ap_arb_share_set_values))) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(cnApi_Av2Av_0_ap_arb_share_counter) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cnApi_Av2Av_0_ap_arb_share_counter))) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))));
  --cnApi_Av2Av_0_ap_allgrants all slave grants, which is an e_mux
  cnApi_Av2Av_0_ap_allgrants <= cnApi_Av2Av_0_ap_grant_vector;
  --cnApi_Av2Av_0_ap_end_xfer assignment, which is an e_assign
  cnApi_Av2Av_0_ap_end_xfer <= NOT ((cnApi_Av2Av_0_ap_waits_for_read OR cnApi_Av2Av_0_ap_waits_for_write));
  --end_xfer_arb_share_counter_term_cnApi_Av2Av_0_ap arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_cnApi_Av2Av_0_ap <= cnApi_Av2Av_0_ap_end_xfer AND (((NOT cnApi_Av2Av_0_ap_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --cnApi_Av2Av_0_ap_arb_share_counter arbitration counter enable, which is an e_assign
  cnApi_Av2Av_0_ap_arb_counter_enable <= ((end_xfer_arb_share_counter_term_cnApi_Av2Av_0_ap AND cnApi_Av2Av_0_ap_allgrants)) OR ((end_xfer_arb_share_counter_term_cnApi_Av2Av_0_ap AND NOT cnApi_Av2Av_0_ap_non_bursting_master_requests));
  --cnApi_Av2Av_0_ap_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      cnApi_Av2Av_0_ap_arb_share_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(cnApi_Av2Av_0_ap_arb_counter_enable) = '1' then 
        cnApi_Av2Av_0_ap_arb_share_counter <= cnApi_Av2Av_0_ap_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --cnApi_Av2Av_0_ap_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      cnApi_Av2Av_0_ap_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((cnApi_Av2Av_0_ap_master_qreq_vector AND end_xfer_arb_share_counter_term_cnApi_Av2Av_0_ap)) OR ((end_xfer_arb_share_counter_term_cnApi_Av2Av_0_ap AND NOT cnApi_Av2Av_0_ap_non_bursting_master_requests)))) = '1' then 
        cnApi_Av2Av_0_ap_slavearbiterlockenable <= cnApi_Av2Av_0_ap_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --ap_cpu/data_master cnApi_Av2Av_0/ap arbiterlock, which is an e_assign
  ap_cpu_data_master_arbiterlock <= cnApi_Av2Av_0_ap_slavearbiterlockenable AND ap_cpu_data_master_continuerequest;
  --cnApi_Av2Av_0_ap_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  cnApi_Av2Av_0_ap_slavearbiterlockenable2 <= cnApi_Av2Av_0_ap_arb_share_counter_next_value;
  --ap_cpu/data_master cnApi_Av2Av_0/ap arbiterlock2, which is an e_assign
  ap_cpu_data_master_arbiterlock2 <= cnApi_Av2Av_0_ap_slavearbiterlockenable2 AND ap_cpu_data_master_continuerequest;
  --cnApi_Av2Av_0_ap_any_continuerequest at least one master continues requesting, which is an e_assign
  cnApi_Av2Av_0_ap_any_continuerequest <= std_logic'('1');
  --ap_cpu_data_master_continuerequest continued request, which is an e_assign
  ap_cpu_data_master_continuerequest <= std_logic'('1');
  internal_ap_cpu_data_master_qualified_request_cnApi_Av2Av_0_ap <= internal_ap_cpu_data_master_requests_cnApi_Av2Av_0_ap AND NOT (((NOT ap_cpu_data_master_waitrequest) AND ap_cpu_data_master_write));
  --cnApi_Av2Av_0_ap_writedata mux, which is an e_mux
  cnApi_Av2Av_0_ap_writedata <= ap_cpu_data_master_writedata;
  --master is always granted when requested
  internal_ap_cpu_data_master_granted_cnApi_Av2Av_0_ap <= internal_ap_cpu_data_master_qualified_request_cnApi_Av2Av_0_ap;
  --ap_cpu/data_master saved-grant cnApi_Av2Av_0/ap, which is an e_assign
  ap_cpu_data_master_saved_grant_cnApi_Av2Av_0_ap <= internal_ap_cpu_data_master_requests_cnApi_Av2Av_0_ap;
  --allow new arb cycle for cnApi_Av2Av_0/ap, which is an e_assign
  cnApi_Av2Av_0_ap_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  cnApi_Av2Av_0_ap_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  cnApi_Av2Av_0_ap_master_qreq_vector <= std_logic'('1');
  --~cnApi_Av2Av_0_ap_reset assignment, which is an e_assign
  cnApi_Av2Av_0_ap_reset <= NOT reset_n;
  cnApi_Av2Av_0_ap_chipselect <= internal_ap_cpu_data_master_granted_cnApi_Av2Av_0_ap;
  --cnApi_Av2Av_0_ap_firsttransfer first transaction, which is an e_assign
  cnApi_Av2Av_0_ap_firsttransfer <= A_WE_StdLogic((std_logic'(cnApi_Av2Av_0_ap_begins_xfer) = '1'), cnApi_Av2Av_0_ap_unreg_firsttransfer, cnApi_Av2Av_0_ap_reg_firsttransfer);
  --cnApi_Av2Av_0_ap_unreg_firsttransfer first transaction, which is an e_assign
  cnApi_Av2Av_0_ap_unreg_firsttransfer <= NOT ((cnApi_Av2Av_0_ap_slavearbiterlockenable AND cnApi_Av2Av_0_ap_any_continuerequest));
  --cnApi_Av2Av_0_ap_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      cnApi_Av2Av_0_ap_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(cnApi_Av2Av_0_ap_begins_xfer) = '1' then 
        cnApi_Av2Av_0_ap_reg_firsttransfer <= cnApi_Av2Av_0_ap_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --cnApi_Av2Av_0_ap_beginbursttransfer_internal begin burst transfer, which is an e_assign
  cnApi_Av2Av_0_ap_beginbursttransfer_internal <= cnApi_Av2Av_0_ap_begins_xfer;
  --cnApi_Av2Av_0_ap_read assignment, which is an e_mux
  cnApi_Av2Av_0_ap_read <= internal_ap_cpu_data_master_granted_cnApi_Av2Av_0_ap AND ap_cpu_data_master_read;
  --cnApi_Av2Av_0_ap_write assignment, which is an e_mux
  cnApi_Av2Av_0_ap_write <= internal_ap_cpu_data_master_granted_cnApi_Av2Av_0_ap AND ap_cpu_data_master_write;
  shifted_address_to_cnApi_Av2Av_0_ap_from_ap_cpu_data_master <= ap_cpu_data_master_address_to_slave;
  --cnApi_Av2Av_0_ap_address mux, which is an e_mux
  cnApi_Av2Av_0_ap_address <= A_EXT (A_SRL(shifted_address_to_cnApi_Av2Av_0_ap_from_ap_cpu_data_master,std_logic_vector'("00000000000000000000000000000010")), 15);
  --d1_cnApi_Av2Av_0_ap_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_cnApi_Av2Av_0_ap_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_cnApi_Av2Av_0_ap_end_xfer <= cnApi_Av2Av_0_ap_end_xfer;
    end if;

  end process;

  --cnApi_Av2Av_0_ap_waits_for_read in a cycle, which is an e_mux
  cnApi_Av2Av_0_ap_waits_for_read <= cnApi_Av2Av_0_ap_in_a_read_cycle AND wait_for_cnApi_Av2Av_0_ap_counter;
  --cnApi_Av2Av_0_ap_in_a_read_cycle assignment, which is an e_assign
  cnApi_Av2Av_0_ap_in_a_read_cycle <= internal_ap_cpu_data_master_granted_cnApi_Av2Av_0_ap AND ap_cpu_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= cnApi_Av2Av_0_ap_in_a_read_cycle;
  --cnApi_Av2Av_0_ap_waits_for_write in a cycle, which is an e_mux
  cnApi_Av2Av_0_ap_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cnApi_Av2Av_0_ap_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --cnApi_Av2Av_0_ap_in_a_write_cycle assignment, which is an e_assign
  cnApi_Av2Av_0_ap_in_a_write_cycle <= internal_ap_cpu_data_master_granted_cnApi_Av2Av_0_ap AND ap_cpu_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= cnApi_Av2Av_0_ap_in_a_write_cycle;
  internal_cnApi_Av2Av_0_ap_wait_counter_eq_0 <= to_std_logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cnApi_Av2Av_0_ap_wait_counter))) = std_logic_vector'("00000000000000000000000000000000")));
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      cnApi_Av2Av_0_ap_wait_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      cnApi_Av2Av_0_ap_wait_counter <= cnApi_Av2Av_0_ap_counter_load_value;
    end if;

  end process;

  cnApi_Av2Av_0_ap_counter_load_value <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(((cnApi_Av2Av_0_ap_in_a_read_cycle AND cnApi_Av2Av_0_ap_begins_xfer))) = '1'), std_logic_vector'("000000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'((NOT internal_cnApi_Av2Av_0_ap_wait_counter_eq_0)) = '1'), ((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cnApi_Av2Av_0_ap_wait_counter))) - std_logic_vector'("000000000000000000000000000000001")), std_logic_vector'("000000000000000000000000000000000"))));
  wait_for_cnApi_Av2Av_0_ap_counter <= cnApi_Av2Av_0_ap_begins_xfer OR NOT internal_cnApi_Av2Av_0_ap_wait_counter_eq_0;
  --cnApi_Av2Av_0_ap_byteenable byte enable port mux, which is an e_mux
  cnApi_Av2Av_0_ap_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_ap_cpu_data_master_granted_cnApi_Av2Av_0_ap)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (ap_cpu_data_master_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))), 4);
  --vhdl renameroo for output signals
  ap_cpu_data_master_granted_cnApi_Av2Av_0_ap <= internal_ap_cpu_data_master_granted_cnApi_Av2Av_0_ap;
  --vhdl renameroo for output signals
  ap_cpu_data_master_qualified_request_cnApi_Av2Av_0_ap <= internal_ap_cpu_data_master_qualified_request_cnApi_Av2Av_0_ap;
  --vhdl renameroo for output signals
  ap_cpu_data_master_requests_cnApi_Av2Av_0_ap <= internal_ap_cpu_data_master_requests_cnApi_Av2Av_0_ap;
  --vhdl renameroo for output signals
  cnApi_Av2Av_0_ap_wait_counter_eq_0 <= internal_cnApi_Av2Av_0_ap_wait_counter_eq_0;
--synthesis translate_off
    --cnApi_Av2Av_0/ap enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity cnApi_Av2Av_0_pcp_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cnApi_Av2Av_0_pcp_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal pcp_cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (25 DOWNTO 0);
                 signal pcp_cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal pcp_cpu_data_master_read : IN STD_LOGIC;
                 signal pcp_cpu_data_master_waitrequest : IN STD_LOGIC;
                 signal pcp_cpu_data_master_write : IN STD_LOGIC;
                 signal pcp_cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cnApi_Av2Av_0_pcp_address : OUT STD_LOGIC_VECTOR (14 DOWNTO 0);
                 signal cnApi_Av2Av_0_pcp_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cnApi_Av2Av_0_pcp_chipselect : OUT STD_LOGIC;
                 signal cnApi_Av2Av_0_pcp_read : OUT STD_LOGIC;
                 signal cnApi_Av2Av_0_pcp_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal cnApi_Av2Av_0_pcp_reset : OUT STD_LOGIC;
                 signal cnApi_Av2Av_0_pcp_wait_counter_eq_0 : OUT STD_LOGIC;
                 signal cnApi_Av2Av_0_pcp_write : OUT STD_LOGIC;
                 signal cnApi_Av2Av_0_pcp_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal d1_cnApi_Av2Av_0_pcp_end_xfer : OUT STD_LOGIC;
                 signal pcp_cpu_data_master_granted_cnApi_Av2Av_0_pcp : OUT STD_LOGIC;
                 signal pcp_cpu_data_master_qualified_request_cnApi_Av2Av_0_pcp : OUT STD_LOGIC;
                 signal pcp_cpu_data_master_read_data_valid_cnApi_Av2Av_0_pcp : OUT STD_LOGIC;
                 signal pcp_cpu_data_master_requests_cnApi_Av2Av_0_pcp : OUT STD_LOGIC
              );
end entity cnApi_Av2Av_0_pcp_arbitrator;


architecture europa of cnApi_Av2Av_0_pcp_arbitrator is
                signal cnApi_Av2Av_0_pcp_allgrants :  STD_LOGIC;
                signal cnApi_Av2Av_0_pcp_allow_new_arb_cycle :  STD_LOGIC;
                signal cnApi_Av2Av_0_pcp_any_bursting_master_saved_grant :  STD_LOGIC;
                signal cnApi_Av2Av_0_pcp_any_continuerequest :  STD_LOGIC;
                signal cnApi_Av2Av_0_pcp_arb_counter_enable :  STD_LOGIC;
                signal cnApi_Av2Av_0_pcp_arb_share_counter :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal cnApi_Av2Av_0_pcp_arb_share_counter_next_value :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal cnApi_Av2Av_0_pcp_arb_share_set_values :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal cnApi_Av2Av_0_pcp_beginbursttransfer_internal :  STD_LOGIC;
                signal cnApi_Av2Av_0_pcp_begins_xfer :  STD_LOGIC;
                signal cnApi_Av2Av_0_pcp_counter_load_value :  STD_LOGIC;
                signal cnApi_Av2Av_0_pcp_end_xfer :  STD_LOGIC;
                signal cnApi_Av2Av_0_pcp_firsttransfer :  STD_LOGIC;
                signal cnApi_Av2Av_0_pcp_grant_vector :  STD_LOGIC;
                signal cnApi_Av2Av_0_pcp_in_a_read_cycle :  STD_LOGIC;
                signal cnApi_Av2Av_0_pcp_in_a_write_cycle :  STD_LOGIC;
                signal cnApi_Av2Av_0_pcp_master_qreq_vector :  STD_LOGIC;
                signal cnApi_Av2Av_0_pcp_non_bursting_master_requests :  STD_LOGIC;
                signal cnApi_Av2Av_0_pcp_reg_firsttransfer :  STD_LOGIC;
                signal cnApi_Av2Av_0_pcp_slavearbiterlockenable :  STD_LOGIC;
                signal cnApi_Av2Av_0_pcp_slavearbiterlockenable2 :  STD_LOGIC;
                signal cnApi_Av2Av_0_pcp_unreg_firsttransfer :  STD_LOGIC;
                signal cnApi_Av2Av_0_pcp_wait_counter :  STD_LOGIC;
                signal cnApi_Av2Av_0_pcp_waits_for_read :  STD_LOGIC;
                signal cnApi_Av2Av_0_pcp_waits_for_write :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_cnApi_Av2Av_0_pcp :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cnApi_Av2Av_0_pcp_wait_counter_eq_0 :  STD_LOGIC;
                signal internal_pcp_cpu_data_master_granted_cnApi_Av2Av_0_pcp :  STD_LOGIC;
                signal internal_pcp_cpu_data_master_qualified_request_cnApi_Av2Av_0_pcp :  STD_LOGIC;
                signal internal_pcp_cpu_data_master_requests_cnApi_Av2Av_0_pcp :  STD_LOGIC;
                signal pcp_cpu_data_master_arbiterlock :  STD_LOGIC;
                signal pcp_cpu_data_master_arbiterlock2 :  STD_LOGIC;
                signal pcp_cpu_data_master_continuerequest :  STD_LOGIC;
                signal pcp_cpu_data_master_saved_grant_cnApi_Av2Av_0_pcp :  STD_LOGIC;
                signal shifted_address_to_cnApi_Av2Av_0_pcp_from_pcp_cpu_data_master :  STD_LOGIC_VECTOR (25 DOWNTO 0);
                signal wait_for_cnApi_Av2Av_0_pcp_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT cnApi_Av2Av_0_pcp_end_xfer;
    end if;

  end process;

  cnApi_Av2Av_0_pcp_begins_xfer <= NOT d1_reasons_to_wait AND (internal_pcp_cpu_data_master_qualified_request_cnApi_Av2Av_0_pcp);
  --assign cnApi_Av2Av_0_pcp_readdata_from_sa = cnApi_Av2Av_0_pcp_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  cnApi_Av2Av_0_pcp_readdata_from_sa <= cnApi_Av2Av_0_pcp_readdata;
  internal_pcp_cpu_data_master_requests_cnApi_Av2Av_0_pcp <= to_std_logic(((Std_Logic_Vector'(pcp_cpu_data_master_address_to_slave(25 DOWNTO 17) & std_logic_vector'("00000000000000000")) = std_logic_vector'("00000000100000000000000000")))) AND ((pcp_cpu_data_master_read OR pcp_cpu_data_master_write));
  --cnApi_Av2Av_0_pcp_arb_share_counter set values, which is an e_mux
  cnApi_Av2Av_0_pcp_arb_share_set_values <= std_logic_vector'("01");
  --cnApi_Av2Av_0_pcp_non_bursting_master_requests mux, which is an e_mux
  cnApi_Av2Av_0_pcp_non_bursting_master_requests <= internal_pcp_cpu_data_master_requests_cnApi_Av2Av_0_pcp;
  --cnApi_Av2Av_0_pcp_any_bursting_master_saved_grant mux, which is an e_mux
  cnApi_Av2Av_0_pcp_any_bursting_master_saved_grant <= std_logic'('0');
  --cnApi_Av2Av_0_pcp_arb_share_counter_next_value assignment, which is an e_assign
  cnApi_Av2Av_0_pcp_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(cnApi_Av2Av_0_pcp_firsttransfer) = '1'), (((std_logic_vector'("0000000000000000000000000000000") & (cnApi_Av2Av_0_pcp_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(cnApi_Av2Av_0_pcp_arb_share_counter)) = '1'), (((std_logic_vector'("0000000000000000000000000000000") & (cnApi_Av2Av_0_pcp_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 2);
  --cnApi_Av2Av_0_pcp_allgrants all slave grants, which is an e_mux
  cnApi_Av2Av_0_pcp_allgrants <= cnApi_Av2Av_0_pcp_grant_vector;
  --cnApi_Av2Av_0_pcp_end_xfer assignment, which is an e_assign
  cnApi_Av2Av_0_pcp_end_xfer <= NOT ((cnApi_Av2Av_0_pcp_waits_for_read OR cnApi_Av2Av_0_pcp_waits_for_write));
  --end_xfer_arb_share_counter_term_cnApi_Av2Av_0_pcp arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_cnApi_Av2Av_0_pcp <= cnApi_Av2Av_0_pcp_end_xfer AND (((NOT cnApi_Av2Av_0_pcp_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --cnApi_Av2Av_0_pcp_arb_share_counter arbitration counter enable, which is an e_assign
  cnApi_Av2Av_0_pcp_arb_counter_enable <= ((end_xfer_arb_share_counter_term_cnApi_Av2Av_0_pcp AND cnApi_Av2Av_0_pcp_allgrants)) OR ((end_xfer_arb_share_counter_term_cnApi_Av2Av_0_pcp AND NOT cnApi_Av2Av_0_pcp_non_bursting_master_requests));
  --cnApi_Av2Av_0_pcp_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      cnApi_Av2Av_0_pcp_arb_share_counter <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      if std_logic'(cnApi_Av2Av_0_pcp_arb_counter_enable) = '1' then 
        cnApi_Av2Av_0_pcp_arb_share_counter <= cnApi_Av2Av_0_pcp_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --cnApi_Av2Av_0_pcp_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      cnApi_Av2Av_0_pcp_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((cnApi_Av2Av_0_pcp_master_qreq_vector AND end_xfer_arb_share_counter_term_cnApi_Av2Av_0_pcp)) OR ((end_xfer_arb_share_counter_term_cnApi_Av2Av_0_pcp AND NOT cnApi_Av2Av_0_pcp_non_bursting_master_requests)))) = '1' then 
        cnApi_Av2Av_0_pcp_slavearbiterlockenable <= or_reduce(cnApi_Av2Av_0_pcp_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --pcp_cpu/data_master cnApi_Av2Av_0/pcp arbiterlock, which is an e_assign
  pcp_cpu_data_master_arbiterlock <= cnApi_Av2Av_0_pcp_slavearbiterlockenable AND pcp_cpu_data_master_continuerequest;
  --cnApi_Av2Av_0_pcp_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  cnApi_Av2Av_0_pcp_slavearbiterlockenable2 <= or_reduce(cnApi_Av2Av_0_pcp_arb_share_counter_next_value);
  --pcp_cpu/data_master cnApi_Av2Av_0/pcp arbiterlock2, which is an e_assign
  pcp_cpu_data_master_arbiterlock2 <= cnApi_Av2Av_0_pcp_slavearbiterlockenable2 AND pcp_cpu_data_master_continuerequest;
  --cnApi_Av2Av_0_pcp_any_continuerequest at least one master continues requesting, which is an e_assign
  cnApi_Av2Av_0_pcp_any_continuerequest <= std_logic'('1');
  --pcp_cpu_data_master_continuerequest continued request, which is an e_assign
  pcp_cpu_data_master_continuerequest <= std_logic'('1');
  internal_pcp_cpu_data_master_qualified_request_cnApi_Av2Av_0_pcp <= internal_pcp_cpu_data_master_requests_cnApi_Av2Av_0_pcp AND NOT (((NOT pcp_cpu_data_master_waitrequest) AND pcp_cpu_data_master_write));
  --cnApi_Av2Av_0_pcp_writedata mux, which is an e_mux
  cnApi_Av2Av_0_pcp_writedata <= pcp_cpu_data_master_writedata;
  --master is always granted when requested
  internal_pcp_cpu_data_master_granted_cnApi_Av2Av_0_pcp <= internal_pcp_cpu_data_master_qualified_request_cnApi_Av2Av_0_pcp;
  --pcp_cpu/data_master saved-grant cnApi_Av2Av_0/pcp, which is an e_assign
  pcp_cpu_data_master_saved_grant_cnApi_Av2Av_0_pcp <= internal_pcp_cpu_data_master_requests_cnApi_Av2Av_0_pcp;
  --allow new arb cycle for cnApi_Av2Av_0/pcp, which is an e_assign
  cnApi_Av2Av_0_pcp_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  cnApi_Av2Av_0_pcp_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  cnApi_Av2Av_0_pcp_master_qreq_vector <= std_logic'('1');
  --~cnApi_Av2Av_0_pcp_reset assignment, which is an e_assign
  cnApi_Av2Av_0_pcp_reset <= NOT reset_n;
  cnApi_Av2Av_0_pcp_chipselect <= internal_pcp_cpu_data_master_granted_cnApi_Av2Av_0_pcp;
  --cnApi_Av2Av_0_pcp_firsttransfer first transaction, which is an e_assign
  cnApi_Av2Av_0_pcp_firsttransfer <= A_WE_StdLogic((std_logic'(cnApi_Av2Av_0_pcp_begins_xfer) = '1'), cnApi_Av2Av_0_pcp_unreg_firsttransfer, cnApi_Av2Av_0_pcp_reg_firsttransfer);
  --cnApi_Av2Av_0_pcp_unreg_firsttransfer first transaction, which is an e_assign
  cnApi_Av2Av_0_pcp_unreg_firsttransfer <= NOT ((cnApi_Av2Av_0_pcp_slavearbiterlockenable AND cnApi_Av2Av_0_pcp_any_continuerequest));
  --cnApi_Av2Av_0_pcp_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      cnApi_Av2Av_0_pcp_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(cnApi_Av2Av_0_pcp_begins_xfer) = '1' then 
        cnApi_Av2Av_0_pcp_reg_firsttransfer <= cnApi_Av2Av_0_pcp_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --cnApi_Av2Av_0_pcp_beginbursttransfer_internal begin burst transfer, which is an e_assign
  cnApi_Av2Av_0_pcp_beginbursttransfer_internal <= cnApi_Av2Av_0_pcp_begins_xfer;
  --cnApi_Av2Av_0_pcp_read assignment, which is an e_mux
  cnApi_Av2Av_0_pcp_read <= internal_pcp_cpu_data_master_granted_cnApi_Av2Av_0_pcp AND pcp_cpu_data_master_read;
  --cnApi_Av2Av_0_pcp_write assignment, which is an e_mux
  cnApi_Av2Av_0_pcp_write <= internal_pcp_cpu_data_master_granted_cnApi_Av2Av_0_pcp AND pcp_cpu_data_master_write;
  shifted_address_to_cnApi_Av2Av_0_pcp_from_pcp_cpu_data_master <= pcp_cpu_data_master_address_to_slave;
  --cnApi_Av2Av_0_pcp_address mux, which is an e_mux
  cnApi_Av2Av_0_pcp_address <= A_EXT (A_SRL(shifted_address_to_cnApi_Av2Av_0_pcp_from_pcp_cpu_data_master,std_logic_vector'("00000000000000000000000000000010")), 15);
  --d1_cnApi_Av2Av_0_pcp_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_cnApi_Av2Av_0_pcp_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_cnApi_Av2Av_0_pcp_end_xfer <= cnApi_Av2Av_0_pcp_end_xfer;
    end if;

  end process;

  --cnApi_Av2Av_0_pcp_waits_for_read in a cycle, which is an e_mux
  cnApi_Av2Av_0_pcp_waits_for_read <= cnApi_Av2Av_0_pcp_in_a_read_cycle AND wait_for_cnApi_Av2Av_0_pcp_counter;
  --cnApi_Av2Av_0_pcp_in_a_read_cycle assignment, which is an e_assign
  cnApi_Av2Av_0_pcp_in_a_read_cycle <= internal_pcp_cpu_data_master_granted_cnApi_Av2Av_0_pcp AND pcp_cpu_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= cnApi_Av2Av_0_pcp_in_a_read_cycle;
  --cnApi_Av2Av_0_pcp_waits_for_write in a cycle, which is an e_mux
  cnApi_Av2Av_0_pcp_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cnApi_Av2Av_0_pcp_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --cnApi_Av2Av_0_pcp_in_a_write_cycle assignment, which is an e_assign
  cnApi_Av2Av_0_pcp_in_a_write_cycle <= internal_pcp_cpu_data_master_granted_cnApi_Av2Av_0_pcp AND pcp_cpu_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= cnApi_Av2Av_0_pcp_in_a_write_cycle;
  internal_cnApi_Av2Av_0_pcp_wait_counter_eq_0 <= to_std_logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cnApi_Av2Av_0_pcp_wait_counter))) = std_logic_vector'("00000000000000000000000000000000")));
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      cnApi_Av2Av_0_pcp_wait_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      cnApi_Av2Av_0_pcp_wait_counter <= cnApi_Av2Av_0_pcp_counter_load_value;
    end if;

  end process;

  cnApi_Av2Av_0_pcp_counter_load_value <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(((cnApi_Av2Av_0_pcp_in_a_read_cycle AND cnApi_Av2Av_0_pcp_begins_xfer))) = '1'), std_logic_vector'("000000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'((NOT internal_cnApi_Av2Av_0_pcp_wait_counter_eq_0)) = '1'), ((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cnApi_Av2Av_0_pcp_wait_counter))) - std_logic_vector'("000000000000000000000000000000001")), std_logic_vector'("000000000000000000000000000000000"))));
  wait_for_cnApi_Av2Av_0_pcp_counter <= cnApi_Av2Av_0_pcp_begins_xfer OR NOT internal_cnApi_Av2Av_0_pcp_wait_counter_eq_0;
  --cnApi_Av2Av_0_pcp_byteenable byte enable port mux, which is an e_mux
  cnApi_Av2Av_0_pcp_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_pcp_cpu_data_master_granted_cnApi_Av2Av_0_pcp)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (pcp_cpu_data_master_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))), 4);
  --vhdl renameroo for output signals
  cnApi_Av2Av_0_pcp_wait_counter_eq_0 <= internal_cnApi_Av2Av_0_pcp_wait_counter_eq_0;
  --vhdl renameroo for output signals
  pcp_cpu_data_master_granted_cnApi_Av2Av_0_pcp <= internal_pcp_cpu_data_master_granted_cnApi_Av2Av_0_pcp;
  --vhdl renameroo for output signals
  pcp_cpu_data_master_qualified_request_cnApi_Av2Av_0_pcp <= internal_pcp_cpu_data_master_qualified_request_cnApi_Av2Av_0_pcp;
  --vhdl renameroo for output signals
  pcp_cpu_data_master_requests_cnApi_Av2Av_0_pcp <= internal_pcp_cpu_data_master_requests_cnApi_Av2Av_0_pcp;
--synthesis translate_off
    --cnApi_Av2Av_0/pcp enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity digio_pio_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal clock_crossing_1_m1_address_to_slave : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal clock_crossing_1_m1_latency_counter : IN STD_LOGIC;
                 signal clock_crossing_1_m1_nativeaddress : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
                 signal clock_crossing_1_m1_read : IN STD_LOGIC;
                 signal clock_crossing_1_m1_write : IN STD_LOGIC;
                 signal clock_crossing_1_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal digio_pio_s1_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal clock_crossing_1_m1_granted_digio_pio_s1 : OUT STD_LOGIC;
                 signal clock_crossing_1_m1_qualified_request_digio_pio_s1 : OUT STD_LOGIC;
                 signal clock_crossing_1_m1_read_data_valid_digio_pio_s1 : OUT STD_LOGIC;
                 signal clock_crossing_1_m1_requests_digio_pio_s1 : OUT STD_LOGIC;
                 signal d1_digio_pio_s1_end_xfer : OUT STD_LOGIC;
                 signal digio_pio_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal digio_pio_s1_chipselect : OUT STD_LOGIC;
                 signal digio_pio_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal digio_pio_s1_reset_n : OUT STD_LOGIC;
                 signal digio_pio_s1_write_n : OUT STD_LOGIC;
                 signal digio_pio_s1_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
              );
end entity digio_pio_s1_arbitrator;


architecture europa of digio_pio_s1_arbitrator is
                signal clock_crossing_1_m1_arbiterlock :  STD_LOGIC;
                signal clock_crossing_1_m1_arbiterlock2 :  STD_LOGIC;
                signal clock_crossing_1_m1_continuerequest :  STD_LOGIC;
                signal clock_crossing_1_m1_saved_grant_digio_pio_s1 :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal digio_pio_s1_allgrants :  STD_LOGIC;
                signal digio_pio_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal digio_pio_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal digio_pio_s1_any_continuerequest :  STD_LOGIC;
                signal digio_pio_s1_arb_counter_enable :  STD_LOGIC;
                signal digio_pio_s1_arb_share_counter :  STD_LOGIC;
                signal digio_pio_s1_arb_share_counter_next_value :  STD_LOGIC;
                signal digio_pio_s1_arb_share_set_values :  STD_LOGIC;
                signal digio_pio_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal digio_pio_s1_begins_xfer :  STD_LOGIC;
                signal digio_pio_s1_end_xfer :  STD_LOGIC;
                signal digio_pio_s1_firsttransfer :  STD_LOGIC;
                signal digio_pio_s1_grant_vector :  STD_LOGIC;
                signal digio_pio_s1_in_a_read_cycle :  STD_LOGIC;
                signal digio_pio_s1_in_a_write_cycle :  STD_LOGIC;
                signal digio_pio_s1_master_qreq_vector :  STD_LOGIC;
                signal digio_pio_s1_non_bursting_master_requests :  STD_LOGIC;
                signal digio_pio_s1_reg_firsttransfer :  STD_LOGIC;
                signal digio_pio_s1_slavearbiterlockenable :  STD_LOGIC;
                signal digio_pio_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal digio_pio_s1_unreg_firsttransfer :  STD_LOGIC;
                signal digio_pio_s1_waits_for_read :  STD_LOGIC;
                signal digio_pio_s1_waits_for_write :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_digio_pio_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_clock_crossing_1_m1_granted_digio_pio_s1 :  STD_LOGIC;
                signal internal_clock_crossing_1_m1_qualified_request_digio_pio_s1 :  STD_LOGIC;
                signal internal_clock_crossing_1_m1_requests_digio_pio_s1 :  STD_LOGIC;
                signal wait_for_digio_pio_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT digio_pio_s1_end_xfer;
    end if;

  end process;

  digio_pio_s1_begins_xfer <= NOT d1_reasons_to_wait AND (internal_clock_crossing_1_m1_qualified_request_digio_pio_s1);
  --assign digio_pio_s1_readdata_from_sa = digio_pio_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  digio_pio_s1_readdata_from_sa <= digio_pio_s1_readdata;
  internal_clock_crossing_1_m1_requests_digio_pio_s1 <= to_std_logic(((Std_Logic_Vector'(clock_crossing_1_m1_address_to_slave(7 DOWNTO 4) & std_logic_vector'("0000")) = std_logic_vector'("10100000")))) AND ((clock_crossing_1_m1_read OR clock_crossing_1_m1_write));
  --digio_pio_s1_arb_share_counter set values, which is an e_mux
  digio_pio_s1_arb_share_set_values <= std_logic'('1');
  --digio_pio_s1_non_bursting_master_requests mux, which is an e_mux
  digio_pio_s1_non_bursting_master_requests <= internal_clock_crossing_1_m1_requests_digio_pio_s1;
  --digio_pio_s1_any_bursting_master_saved_grant mux, which is an e_mux
  digio_pio_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --digio_pio_s1_arb_share_counter_next_value assignment, which is an e_assign
  digio_pio_s1_arb_share_counter_next_value <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(digio_pio_s1_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(digio_pio_s1_arb_share_set_values))) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(digio_pio_s1_arb_share_counter) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(digio_pio_s1_arb_share_counter))) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))));
  --digio_pio_s1_allgrants all slave grants, which is an e_mux
  digio_pio_s1_allgrants <= digio_pio_s1_grant_vector;
  --digio_pio_s1_end_xfer assignment, which is an e_assign
  digio_pio_s1_end_xfer <= NOT ((digio_pio_s1_waits_for_read OR digio_pio_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_digio_pio_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_digio_pio_s1 <= digio_pio_s1_end_xfer AND (((NOT digio_pio_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --digio_pio_s1_arb_share_counter arbitration counter enable, which is an e_assign
  digio_pio_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_digio_pio_s1 AND digio_pio_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_digio_pio_s1 AND NOT digio_pio_s1_non_bursting_master_requests));
  --digio_pio_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      digio_pio_s1_arb_share_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(digio_pio_s1_arb_counter_enable) = '1' then 
        digio_pio_s1_arb_share_counter <= digio_pio_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --digio_pio_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      digio_pio_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((digio_pio_s1_master_qreq_vector AND end_xfer_arb_share_counter_term_digio_pio_s1)) OR ((end_xfer_arb_share_counter_term_digio_pio_s1 AND NOT digio_pio_s1_non_bursting_master_requests)))) = '1' then 
        digio_pio_s1_slavearbiterlockenable <= digio_pio_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --clock_crossing_1/m1 digio_pio/s1 arbiterlock, which is an e_assign
  clock_crossing_1_m1_arbiterlock <= digio_pio_s1_slavearbiterlockenable AND clock_crossing_1_m1_continuerequest;
  --digio_pio_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  digio_pio_s1_slavearbiterlockenable2 <= digio_pio_s1_arb_share_counter_next_value;
  --clock_crossing_1/m1 digio_pio/s1 arbiterlock2, which is an e_assign
  clock_crossing_1_m1_arbiterlock2 <= digio_pio_s1_slavearbiterlockenable2 AND clock_crossing_1_m1_continuerequest;
  --digio_pio_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  digio_pio_s1_any_continuerequest <= std_logic'('1');
  --clock_crossing_1_m1_continuerequest continued request, which is an e_assign
  clock_crossing_1_m1_continuerequest <= std_logic'('1');
  internal_clock_crossing_1_m1_qualified_request_digio_pio_s1 <= internal_clock_crossing_1_m1_requests_digio_pio_s1 AND NOT ((clock_crossing_1_m1_read AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(clock_crossing_1_m1_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))))));
  --local readdatavalid clock_crossing_1_m1_read_data_valid_digio_pio_s1, which is an e_mux
  clock_crossing_1_m1_read_data_valid_digio_pio_s1 <= (internal_clock_crossing_1_m1_granted_digio_pio_s1 AND clock_crossing_1_m1_read) AND NOT digio_pio_s1_waits_for_read;
  --digio_pio_s1_writedata mux, which is an e_mux
  digio_pio_s1_writedata <= clock_crossing_1_m1_writedata;
  --master is always granted when requested
  internal_clock_crossing_1_m1_granted_digio_pio_s1 <= internal_clock_crossing_1_m1_qualified_request_digio_pio_s1;
  --clock_crossing_1/m1 saved-grant digio_pio/s1, which is an e_assign
  clock_crossing_1_m1_saved_grant_digio_pio_s1 <= internal_clock_crossing_1_m1_requests_digio_pio_s1;
  --allow new arb cycle for digio_pio/s1, which is an e_assign
  digio_pio_s1_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  digio_pio_s1_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  digio_pio_s1_master_qreq_vector <= std_logic'('1');
  --digio_pio_s1_reset_n assignment, which is an e_assign
  digio_pio_s1_reset_n <= reset_n;
  digio_pio_s1_chipselect <= internal_clock_crossing_1_m1_granted_digio_pio_s1;
  --digio_pio_s1_firsttransfer first transaction, which is an e_assign
  digio_pio_s1_firsttransfer <= A_WE_StdLogic((std_logic'(digio_pio_s1_begins_xfer) = '1'), digio_pio_s1_unreg_firsttransfer, digio_pio_s1_reg_firsttransfer);
  --digio_pio_s1_unreg_firsttransfer first transaction, which is an e_assign
  digio_pio_s1_unreg_firsttransfer <= NOT ((digio_pio_s1_slavearbiterlockenable AND digio_pio_s1_any_continuerequest));
  --digio_pio_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      digio_pio_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(digio_pio_s1_begins_xfer) = '1' then 
        digio_pio_s1_reg_firsttransfer <= digio_pio_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --digio_pio_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  digio_pio_s1_beginbursttransfer_internal <= digio_pio_s1_begins_xfer;
  --~digio_pio_s1_write_n assignment, which is an e_mux
  digio_pio_s1_write_n <= NOT ((internal_clock_crossing_1_m1_granted_digio_pio_s1 AND clock_crossing_1_m1_write));
  --digio_pio_s1_address mux, which is an e_mux
  digio_pio_s1_address <= clock_crossing_1_m1_nativeaddress (1 DOWNTO 0);
  --d1_digio_pio_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_digio_pio_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_digio_pio_s1_end_xfer <= digio_pio_s1_end_xfer;
    end if;

  end process;

  --digio_pio_s1_waits_for_read in a cycle, which is an e_mux
  digio_pio_s1_waits_for_read <= digio_pio_s1_in_a_read_cycle AND digio_pio_s1_begins_xfer;
  --digio_pio_s1_in_a_read_cycle assignment, which is an e_assign
  digio_pio_s1_in_a_read_cycle <= internal_clock_crossing_1_m1_granted_digio_pio_s1 AND clock_crossing_1_m1_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= digio_pio_s1_in_a_read_cycle;
  --digio_pio_s1_waits_for_write in a cycle, which is an e_mux
  digio_pio_s1_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(digio_pio_s1_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --digio_pio_s1_in_a_write_cycle assignment, which is an e_assign
  digio_pio_s1_in_a_write_cycle <= internal_clock_crossing_1_m1_granted_digio_pio_s1 AND clock_crossing_1_m1_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= digio_pio_s1_in_a_write_cycle;
  wait_for_digio_pio_s1_counter <= std_logic'('0');
  --vhdl renameroo for output signals
  clock_crossing_1_m1_granted_digio_pio_s1 <= internal_clock_crossing_1_m1_granted_digio_pio_s1;
  --vhdl renameroo for output signals
  clock_crossing_1_m1_qualified_request_digio_pio_s1 <= internal_clock_crossing_1_m1_qualified_request_digio_pio_s1;
  --vhdl renameroo for output signals
  clock_crossing_1_m1_requests_digio_pio_s1 <= internal_clock_crossing_1_m1_requests_digio_pio_s1;
--synthesis translate_off
    --digio_pio/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity epcs_flash_controller_0_epcs_control_port_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal epcs_flash_controller_0_epcs_control_port_dataavailable : IN STD_LOGIC;
                 signal epcs_flash_controller_0_epcs_control_port_endofpacket : IN STD_LOGIC;
                 signal epcs_flash_controller_0_epcs_control_port_irq : IN STD_LOGIC;
                 signal epcs_flash_controller_0_epcs_control_port_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal epcs_flash_controller_0_epcs_control_port_readyfordata : IN STD_LOGIC;
                 signal pcp_cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (25 DOWNTO 0);
                 signal pcp_cpu_data_master_read : IN STD_LOGIC;
                 signal pcp_cpu_data_master_write : IN STD_LOGIC;
                 signal pcp_cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal pcp_cpu_instruction_master_address_to_slave : IN STD_LOGIC_VECTOR (25 DOWNTO 0);
                 signal pcp_cpu_instruction_master_latency_counter : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal pcp_cpu_instruction_master_read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal d1_epcs_flash_controller_0_epcs_control_port_end_xfer : OUT STD_LOGIC;
                 signal epcs_flash_controller_0_epcs_control_port_address : OUT STD_LOGIC_VECTOR (8 DOWNTO 0);
                 signal epcs_flash_controller_0_epcs_control_port_chipselect : OUT STD_LOGIC;
                 signal epcs_flash_controller_0_epcs_control_port_dataavailable_from_sa : OUT STD_LOGIC;
                 signal epcs_flash_controller_0_epcs_control_port_endofpacket_from_sa : OUT STD_LOGIC;
                 signal epcs_flash_controller_0_epcs_control_port_irq_from_sa : OUT STD_LOGIC;
                 signal epcs_flash_controller_0_epcs_control_port_read_n : OUT STD_LOGIC;
                 signal epcs_flash_controller_0_epcs_control_port_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal epcs_flash_controller_0_epcs_control_port_readyfordata_from_sa : OUT STD_LOGIC;
                 signal epcs_flash_controller_0_epcs_control_port_reset_n : OUT STD_LOGIC;
                 signal epcs_flash_controller_0_epcs_control_port_write_n : OUT STD_LOGIC;
                 signal epcs_flash_controller_0_epcs_control_port_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal pcp_cpu_data_master_granted_epcs_flash_controller_0_epcs_control_port : OUT STD_LOGIC;
                 signal pcp_cpu_data_master_qualified_request_epcs_flash_controller_0_epcs_control_port : OUT STD_LOGIC;
                 signal pcp_cpu_data_master_read_data_valid_epcs_flash_controller_0_epcs_control_port : OUT STD_LOGIC;
                 signal pcp_cpu_data_master_requests_epcs_flash_controller_0_epcs_control_port : OUT STD_LOGIC;
                 signal pcp_cpu_instruction_master_granted_epcs_flash_controller_0_epcs_control_port : OUT STD_LOGIC;
                 signal pcp_cpu_instruction_master_qualified_request_epcs_flash_controller_0_epcs_control_port : OUT STD_LOGIC;
                 signal pcp_cpu_instruction_master_read_data_valid_epcs_flash_controller_0_epcs_control_port : OUT STD_LOGIC;
                 signal pcp_cpu_instruction_master_requests_epcs_flash_controller_0_epcs_control_port : OUT STD_LOGIC
              );
end entity epcs_flash_controller_0_epcs_control_port_arbitrator;


architecture europa of epcs_flash_controller_0_epcs_control_port_arbitrator is
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_epcs_flash_controller_0_epcs_control_port :  STD_LOGIC;
                signal epcs_flash_controller_0_epcs_control_port_allgrants :  STD_LOGIC;
                signal epcs_flash_controller_0_epcs_control_port_allow_new_arb_cycle :  STD_LOGIC;
                signal epcs_flash_controller_0_epcs_control_port_any_bursting_master_saved_grant :  STD_LOGIC;
                signal epcs_flash_controller_0_epcs_control_port_any_continuerequest :  STD_LOGIC;
                signal epcs_flash_controller_0_epcs_control_port_arb_addend :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal epcs_flash_controller_0_epcs_control_port_arb_counter_enable :  STD_LOGIC;
                signal epcs_flash_controller_0_epcs_control_port_arb_share_counter :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal epcs_flash_controller_0_epcs_control_port_arb_share_counter_next_value :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal epcs_flash_controller_0_epcs_control_port_arb_share_set_values :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal epcs_flash_controller_0_epcs_control_port_arb_winner :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal epcs_flash_controller_0_epcs_control_port_arbitration_holdoff_internal :  STD_LOGIC;
                signal epcs_flash_controller_0_epcs_control_port_beginbursttransfer_internal :  STD_LOGIC;
                signal epcs_flash_controller_0_epcs_control_port_begins_xfer :  STD_LOGIC;
                signal epcs_flash_controller_0_epcs_control_port_chosen_master_double_vector :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal epcs_flash_controller_0_epcs_control_port_chosen_master_rot_left :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal epcs_flash_controller_0_epcs_control_port_end_xfer :  STD_LOGIC;
                signal epcs_flash_controller_0_epcs_control_port_firsttransfer :  STD_LOGIC;
                signal epcs_flash_controller_0_epcs_control_port_grant_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal epcs_flash_controller_0_epcs_control_port_in_a_read_cycle :  STD_LOGIC;
                signal epcs_flash_controller_0_epcs_control_port_in_a_write_cycle :  STD_LOGIC;
                signal epcs_flash_controller_0_epcs_control_port_master_qreq_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal epcs_flash_controller_0_epcs_control_port_non_bursting_master_requests :  STD_LOGIC;
                signal epcs_flash_controller_0_epcs_control_port_reg_firsttransfer :  STD_LOGIC;
                signal epcs_flash_controller_0_epcs_control_port_saved_chosen_master_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal epcs_flash_controller_0_epcs_control_port_slavearbiterlockenable :  STD_LOGIC;
                signal epcs_flash_controller_0_epcs_control_port_slavearbiterlockenable2 :  STD_LOGIC;
                signal epcs_flash_controller_0_epcs_control_port_unreg_firsttransfer :  STD_LOGIC;
                signal epcs_flash_controller_0_epcs_control_port_waits_for_read :  STD_LOGIC;
                signal epcs_flash_controller_0_epcs_control_port_waits_for_write :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_pcp_cpu_data_master_granted_epcs_flash_controller_0_epcs_control_port :  STD_LOGIC;
                signal internal_pcp_cpu_data_master_qualified_request_epcs_flash_controller_0_epcs_control_port :  STD_LOGIC;
                signal internal_pcp_cpu_data_master_requests_epcs_flash_controller_0_epcs_control_port :  STD_LOGIC;
                signal internal_pcp_cpu_instruction_master_granted_epcs_flash_controller_0_epcs_control_port :  STD_LOGIC;
                signal internal_pcp_cpu_instruction_master_qualified_request_epcs_flash_controller_0_epcs_control_port :  STD_LOGIC;
                signal internal_pcp_cpu_instruction_master_requests_epcs_flash_controller_0_epcs_control_port :  STD_LOGIC;
                signal last_cycle_pcp_cpu_data_master_granted_slave_epcs_flash_controller_0_epcs_control_port :  STD_LOGIC;
                signal last_cycle_pcp_cpu_instruction_master_granted_slave_epcs_flash_controller_0_epcs_control_port :  STD_LOGIC;
                signal pcp_cpu_data_master_arbiterlock :  STD_LOGIC;
                signal pcp_cpu_data_master_arbiterlock2 :  STD_LOGIC;
                signal pcp_cpu_data_master_continuerequest :  STD_LOGIC;
                signal pcp_cpu_data_master_saved_grant_epcs_flash_controller_0_epcs_control_port :  STD_LOGIC;
                signal pcp_cpu_instruction_master_arbiterlock :  STD_LOGIC;
                signal pcp_cpu_instruction_master_arbiterlock2 :  STD_LOGIC;
                signal pcp_cpu_instruction_master_continuerequest :  STD_LOGIC;
                signal pcp_cpu_instruction_master_saved_grant_epcs_flash_controller_0_epcs_control_port :  STD_LOGIC;
                signal shifted_address_to_epcs_flash_controller_0_epcs_control_port_from_pcp_cpu_data_master :  STD_LOGIC_VECTOR (25 DOWNTO 0);
                signal shifted_address_to_epcs_flash_controller_0_epcs_control_port_from_pcp_cpu_instruction_master :  STD_LOGIC_VECTOR (25 DOWNTO 0);
                signal wait_for_epcs_flash_controller_0_epcs_control_port_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT epcs_flash_controller_0_epcs_control_port_end_xfer;
    end if;

  end process;

  epcs_flash_controller_0_epcs_control_port_begins_xfer <= NOT d1_reasons_to_wait AND ((internal_pcp_cpu_data_master_qualified_request_epcs_flash_controller_0_epcs_control_port OR internal_pcp_cpu_instruction_master_qualified_request_epcs_flash_controller_0_epcs_control_port));
  --assign epcs_flash_controller_0_epcs_control_port_readdata_from_sa = epcs_flash_controller_0_epcs_control_port_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  epcs_flash_controller_0_epcs_control_port_readdata_from_sa <= epcs_flash_controller_0_epcs_control_port_readdata;
  internal_pcp_cpu_data_master_requests_epcs_flash_controller_0_epcs_control_port <= to_std_logic(((Std_Logic_Vector'(pcp_cpu_data_master_address_to_slave(25 DOWNTO 11) & std_logic_vector'("00000000000")) = std_logic_vector'("00000000000000000000000000")))) AND ((pcp_cpu_data_master_read OR pcp_cpu_data_master_write));
  --assign epcs_flash_controller_0_epcs_control_port_dataavailable_from_sa = epcs_flash_controller_0_epcs_control_port_dataavailable so that symbol knows where to group signals which may go to master only, which is an e_assign
  epcs_flash_controller_0_epcs_control_port_dataavailable_from_sa <= epcs_flash_controller_0_epcs_control_port_dataavailable;
  --assign epcs_flash_controller_0_epcs_control_port_readyfordata_from_sa = epcs_flash_controller_0_epcs_control_port_readyfordata so that symbol knows where to group signals which may go to master only, which is an e_assign
  epcs_flash_controller_0_epcs_control_port_readyfordata_from_sa <= epcs_flash_controller_0_epcs_control_port_readyfordata;
  --epcs_flash_controller_0_epcs_control_port_arb_share_counter set values, which is an e_mux
  epcs_flash_controller_0_epcs_control_port_arb_share_set_values <= std_logic_vector'("01");
  --epcs_flash_controller_0_epcs_control_port_non_bursting_master_requests mux, which is an e_mux
  epcs_flash_controller_0_epcs_control_port_non_bursting_master_requests <= ((internal_pcp_cpu_data_master_requests_epcs_flash_controller_0_epcs_control_port OR internal_pcp_cpu_instruction_master_requests_epcs_flash_controller_0_epcs_control_port) OR internal_pcp_cpu_data_master_requests_epcs_flash_controller_0_epcs_control_port) OR internal_pcp_cpu_instruction_master_requests_epcs_flash_controller_0_epcs_control_port;
  --epcs_flash_controller_0_epcs_control_port_any_bursting_master_saved_grant mux, which is an e_mux
  epcs_flash_controller_0_epcs_control_port_any_bursting_master_saved_grant <= std_logic'('0');
  --epcs_flash_controller_0_epcs_control_port_arb_share_counter_next_value assignment, which is an e_assign
  epcs_flash_controller_0_epcs_control_port_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(epcs_flash_controller_0_epcs_control_port_firsttransfer) = '1'), (((std_logic_vector'("0000000000000000000000000000000") & (epcs_flash_controller_0_epcs_control_port_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(epcs_flash_controller_0_epcs_control_port_arb_share_counter)) = '1'), (((std_logic_vector'("0000000000000000000000000000000") & (epcs_flash_controller_0_epcs_control_port_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 2);
  --epcs_flash_controller_0_epcs_control_port_allgrants all slave grants, which is an e_mux
  epcs_flash_controller_0_epcs_control_port_allgrants <= (((or_reduce(epcs_flash_controller_0_epcs_control_port_grant_vector)) OR (or_reduce(epcs_flash_controller_0_epcs_control_port_grant_vector))) OR (or_reduce(epcs_flash_controller_0_epcs_control_port_grant_vector))) OR (or_reduce(epcs_flash_controller_0_epcs_control_port_grant_vector));
  --epcs_flash_controller_0_epcs_control_port_end_xfer assignment, which is an e_assign
  epcs_flash_controller_0_epcs_control_port_end_xfer <= NOT ((epcs_flash_controller_0_epcs_control_port_waits_for_read OR epcs_flash_controller_0_epcs_control_port_waits_for_write));
  --end_xfer_arb_share_counter_term_epcs_flash_controller_0_epcs_control_port arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_epcs_flash_controller_0_epcs_control_port <= epcs_flash_controller_0_epcs_control_port_end_xfer AND (((NOT epcs_flash_controller_0_epcs_control_port_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --epcs_flash_controller_0_epcs_control_port_arb_share_counter arbitration counter enable, which is an e_assign
  epcs_flash_controller_0_epcs_control_port_arb_counter_enable <= ((end_xfer_arb_share_counter_term_epcs_flash_controller_0_epcs_control_port AND epcs_flash_controller_0_epcs_control_port_allgrants)) OR ((end_xfer_arb_share_counter_term_epcs_flash_controller_0_epcs_control_port AND NOT epcs_flash_controller_0_epcs_control_port_non_bursting_master_requests));
  --epcs_flash_controller_0_epcs_control_port_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      epcs_flash_controller_0_epcs_control_port_arb_share_counter <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      if std_logic'(epcs_flash_controller_0_epcs_control_port_arb_counter_enable) = '1' then 
        epcs_flash_controller_0_epcs_control_port_arb_share_counter <= epcs_flash_controller_0_epcs_control_port_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --epcs_flash_controller_0_epcs_control_port_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      epcs_flash_controller_0_epcs_control_port_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((or_reduce(epcs_flash_controller_0_epcs_control_port_master_qreq_vector) AND end_xfer_arb_share_counter_term_epcs_flash_controller_0_epcs_control_port)) OR ((end_xfer_arb_share_counter_term_epcs_flash_controller_0_epcs_control_port AND NOT epcs_flash_controller_0_epcs_control_port_non_bursting_master_requests)))) = '1' then 
        epcs_flash_controller_0_epcs_control_port_slavearbiterlockenable <= or_reduce(epcs_flash_controller_0_epcs_control_port_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --pcp_cpu/data_master epcs_flash_controller_0/epcs_control_port arbiterlock, which is an e_assign
  pcp_cpu_data_master_arbiterlock <= epcs_flash_controller_0_epcs_control_port_slavearbiterlockenable AND pcp_cpu_data_master_continuerequest;
  --epcs_flash_controller_0_epcs_control_port_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  epcs_flash_controller_0_epcs_control_port_slavearbiterlockenable2 <= or_reduce(epcs_flash_controller_0_epcs_control_port_arb_share_counter_next_value);
  --pcp_cpu/data_master epcs_flash_controller_0/epcs_control_port arbiterlock2, which is an e_assign
  pcp_cpu_data_master_arbiterlock2 <= epcs_flash_controller_0_epcs_control_port_slavearbiterlockenable2 AND pcp_cpu_data_master_continuerequest;
  --pcp_cpu/instruction_master epcs_flash_controller_0/epcs_control_port arbiterlock, which is an e_assign
  pcp_cpu_instruction_master_arbiterlock <= epcs_flash_controller_0_epcs_control_port_slavearbiterlockenable AND pcp_cpu_instruction_master_continuerequest;
  --pcp_cpu/instruction_master epcs_flash_controller_0/epcs_control_port arbiterlock2, which is an e_assign
  pcp_cpu_instruction_master_arbiterlock2 <= epcs_flash_controller_0_epcs_control_port_slavearbiterlockenable2 AND pcp_cpu_instruction_master_continuerequest;
  --pcp_cpu/instruction_master granted epcs_flash_controller_0/epcs_control_port last time, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      last_cycle_pcp_cpu_instruction_master_granted_slave_epcs_flash_controller_0_epcs_control_port <= std_logic'('0');
    elsif clk'event and clk = '1' then
      last_cycle_pcp_cpu_instruction_master_granted_slave_epcs_flash_controller_0_epcs_control_port <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(pcp_cpu_instruction_master_saved_grant_epcs_flash_controller_0_epcs_control_port) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((epcs_flash_controller_0_epcs_control_port_arbitration_holdoff_internal OR NOT internal_pcp_cpu_instruction_master_requests_epcs_flash_controller_0_epcs_control_port))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_pcp_cpu_instruction_master_granted_slave_epcs_flash_controller_0_epcs_control_port))))));
    end if;

  end process;

  --pcp_cpu_instruction_master_continuerequest continued request, which is an e_mux
  pcp_cpu_instruction_master_continuerequest <= last_cycle_pcp_cpu_instruction_master_granted_slave_epcs_flash_controller_0_epcs_control_port AND internal_pcp_cpu_instruction_master_requests_epcs_flash_controller_0_epcs_control_port;
  --epcs_flash_controller_0_epcs_control_port_any_continuerequest at least one master continues requesting, which is an e_mux
  epcs_flash_controller_0_epcs_control_port_any_continuerequest <= pcp_cpu_instruction_master_continuerequest OR pcp_cpu_data_master_continuerequest;
  internal_pcp_cpu_data_master_qualified_request_epcs_flash_controller_0_epcs_control_port <= internal_pcp_cpu_data_master_requests_epcs_flash_controller_0_epcs_control_port AND NOT (pcp_cpu_instruction_master_arbiterlock);
  --epcs_flash_controller_0_epcs_control_port_writedata mux, which is an e_mux
  epcs_flash_controller_0_epcs_control_port_writedata <= pcp_cpu_data_master_writedata;
  --assign epcs_flash_controller_0_epcs_control_port_endofpacket_from_sa = epcs_flash_controller_0_epcs_control_port_endofpacket so that symbol knows where to group signals which may go to master only, which is an e_assign
  epcs_flash_controller_0_epcs_control_port_endofpacket_from_sa <= epcs_flash_controller_0_epcs_control_port_endofpacket;
  internal_pcp_cpu_instruction_master_requests_epcs_flash_controller_0_epcs_control_port <= ((to_std_logic(((Std_Logic_Vector'(pcp_cpu_instruction_master_address_to_slave(25 DOWNTO 11) & std_logic_vector'("00000000000")) = std_logic_vector'("00000000000000000000000000")))) AND (pcp_cpu_instruction_master_read))) AND pcp_cpu_instruction_master_read;
  --pcp_cpu/data_master granted epcs_flash_controller_0/epcs_control_port last time, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      last_cycle_pcp_cpu_data_master_granted_slave_epcs_flash_controller_0_epcs_control_port <= std_logic'('0');
    elsif clk'event and clk = '1' then
      last_cycle_pcp_cpu_data_master_granted_slave_epcs_flash_controller_0_epcs_control_port <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(pcp_cpu_data_master_saved_grant_epcs_flash_controller_0_epcs_control_port) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((epcs_flash_controller_0_epcs_control_port_arbitration_holdoff_internal OR NOT internal_pcp_cpu_data_master_requests_epcs_flash_controller_0_epcs_control_port))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_pcp_cpu_data_master_granted_slave_epcs_flash_controller_0_epcs_control_port))))));
    end if;

  end process;

  --pcp_cpu_data_master_continuerequest continued request, which is an e_mux
  pcp_cpu_data_master_continuerequest <= last_cycle_pcp_cpu_data_master_granted_slave_epcs_flash_controller_0_epcs_control_port AND internal_pcp_cpu_data_master_requests_epcs_flash_controller_0_epcs_control_port;
  internal_pcp_cpu_instruction_master_qualified_request_epcs_flash_controller_0_epcs_control_port <= internal_pcp_cpu_instruction_master_requests_epcs_flash_controller_0_epcs_control_port AND NOT ((((pcp_cpu_instruction_master_read AND to_std_logic((((std_logic_vector'("000000000000000000000000000000") & (pcp_cpu_instruction_master_latency_counter)) /= std_logic_vector'("00000000000000000000000000000000")))))) OR pcp_cpu_data_master_arbiterlock));
  --local readdatavalid pcp_cpu_instruction_master_read_data_valid_epcs_flash_controller_0_epcs_control_port, which is an e_mux
  pcp_cpu_instruction_master_read_data_valid_epcs_flash_controller_0_epcs_control_port <= (internal_pcp_cpu_instruction_master_granted_epcs_flash_controller_0_epcs_control_port AND pcp_cpu_instruction_master_read) AND NOT epcs_flash_controller_0_epcs_control_port_waits_for_read;
  --allow new arb cycle for epcs_flash_controller_0/epcs_control_port, which is an e_assign
  epcs_flash_controller_0_epcs_control_port_allow_new_arb_cycle <= NOT pcp_cpu_data_master_arbiterlock AND NOT pcp_cpu_instruction_master_arbiterlock;
  --pcp_cpu/instruction_master assignment into master qualified-requests vector for epcs_flash_controller_0/epcs_control_port, which is an e_assign
  epcs_flash_controller_0_epcs_control_port_master_qreq_vector(0) <= internal_pcp_cpu_instruction_master_qualified_request_epcs_flash_controller_0_epcs_control_port;
  --pcp_cpu/instruction_master grant epcs_flash_controller_0/epcs_control_port, which is an e_assign
  internal_pcp_cpu_instruction_master_granted_epcs_flash_controller_0_epcs_control_port <= epcs_flash_controller_0_epcs_control_port_grant_vector(0);
  --pcp_cpu/instruction_master saved-grant epcs_flash_controller_0/epcs_control_port, which is an e_assign
  pcp_cpu_instruction_master_saved_grant_epcs_flash_controller_0_epcs_control_port <= epcs_flash_controller_0_epcs_control_port_arb_winner(0) AND internal_pcp_cpu_instruction_master_requests_epcs_flash_controller_0_epcs_control_port;
  --pcp_cpu/data_master assignment into master qualified-requests vector for epcs_flash_controller_0/epcs_control_port, which is an e_assign
  epcs_flash_controller_0_epcs_control_port_master_qreq_vector(1) <= internal_pcp_cpu_data_master_qualified_request_epcs_flash_controller_0_epcs_control_port;
  --pcp_cpu/data_master grant epcs_flash_controller_0/epcs_control_port, which is an e_assign
  internal_pcp_cpu_data_master_granted_epcs_flash_controller_0_epcs_control_port <= epcs_flash_controller_0_epcs_control_port_grant_vector(1);
  --pcp_cpu/data_master saved-grant epcs_flash_controller_0/epcs_control_port, which is an e_assign
  pcp_cpu_data_master_saved_grant_epcs_flash_controller_0_epcs_control_port <= epcs_flash_controller_0_epcs_control_port_arb_winner(1) AND internal_pcp_cpu_data_master_requests_epcs_flash_controller_0_epcs_control_port;
  --epcs_flash_controller_0/epcs_control_port chosen-master double-vector, which is an e_assign
  epcs_flash_controller_0_epcs_control_port_chosen_master_double_vector <= A_EXT (((std_logic_vector'("0") & ((epcs_flash_controller_0_epcs_control_port_master_qreq_vector & epcs_flash_controller_0_epcs_control_port_master_qreq_vector))) AND (((std_logic_vector'("0") & (Std_Logic_Vector'(NOT epcs_flash_controller_0_epcs_control_port_master_qreq_vector & NOT epcs_flash_controller_0_epcs_control_port_master_qreq_vector))) + (std_logic_vector'("000") & (epcs_flash_controller_0_epcs_control_port_arb_addend))))), 4);
  --stable onehot encoding of arb winner
  epcs_flash_controller_0_epcs_control_port_arb_winner <= A_WE_StdLogicVector((std_logic'(((epcs_flash_controller_0_epcs_control_port_allow_new_arb_cycle AND or_reduce(epcs_flash_controller_0_epcs_control_port_grant_vector)))) = '1'), epcs_flash_controller_0_epcs_control_port_grant_vector, epcs_flash_controller_0_epcs_control_port_saved_chosen_master_vector);
  --saved epcs_flash_controller_0_epcs_control_port_grant_vector, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      epcs_flash_controller_0_epcs_control_port_saved_chosen_master_vector <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      if std_logic'(epcs_flash_controller_0_epcs_control_port_allow_new_arb_cycle) = '1' then 
        epcs_flash_controller_0_epcs_control_port_saved_chosen_master_vector <= A_WE_StdLogicVector((std_logic'(or_reduce(epcs_flash_controller_0_epcs_control_port_grant_vector)) = '1'), epcs_flash_controller_0_epcs_control_port_grant_vector, epcs_flash_controller_0_epcs_control_port_saved_chosen_master_vector);
      end if;
    end if;

  end process;

  --onehot encoding of chosen master
  epcs_flash_controller_0_epcs_control_port_grant_vector <= Std_Logic_Vector'(A_ToStdLogicVector(((epcs_flash_controller_0_epcs_control_port_chosen_master_double_vector(1) OR epcs_flash_controller_0_epcs_control_port_chosen_master_double_vector(3)))) & A_ToStdLogicVector(((epcs_flash_controller_0_epcs_control_port_chosen_master_double_vector(0) OR epcs_flash_controller_0_epcs_control_port_chosen_master_double_vector(2)))));
  --epcs_flash_controller_0/epcs_control_port chosen master rotated left, which is an e_assign
  epcs_flash_controller_0_epcs_control_port_chosen_master_rot_left <= A_EXT (A_WE_StdLogicVector((((A_SLL(epcs_flash_controller_0_epcs_control_port_arb_winner,std_logic_vector'("00000000000000000000000000000001")))) /= std_logic_vector'("00")), (std_logic_vector'("000000000000000000000000000000") & ((A_SLL(epcs_flash_controller_0_epcs_control_port_arb_winner,std_logic_vector'("00000000000000000000000000000001"))))), std_logic_vector'("00000000000000000000000000000001")), 2);
  --epcs_flash_controller_0/epcs_control_port's addend for next-master-grant
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      epcs_flash_controller_0_epcs_control_port_arb_addend <= std_logic_vector'("01");
    elsif clk'event and clk = '1' then
      if std_logic'(or_reduce(epcs_flash_controller_0_epcs_control_port_grant_vector)) = '1' then 
        epcs_flash_controller_0_epcs_control_port_arb_addend <= A_WE_StdLogicVector((std_logic'(epcs_flash_controller_0_epcs_control_port_end_xfer) = '1'), epcs_flash_controller_0_epcs_control_port_chosen_master_rot_left, epcs_flash_controller_0_epcs_control_port_grant_vector);
      end if;
    end if;

  end process;

  --epcs_flash_controller_0_epcs_control_port_reset_n assignment, which is an e_assign
  epcs_flash_controller_0_epcs_control_port_reset_n <= reset_n;
  epcs_flash_controller_0_epcs_control_port_chipselect <= internal_pcp_cpu_data_master_granted_epcs_flash_controller_0_epcs_control_port OR internal_pcp_cpu_instruction_master_granted_epcs_flash_controller_0_epcs_control_port;
  --epcs_flash_controller_0_epcs_control_port_firsttransfer first transaction, which is an e_assign
  epcs_flash_controller_0_epcs_control_port_firsttransfer <= A_WE_StdLogic((std_logic'(epcs_flash_controller_0_epcs_control_port_begins_xfer) = '1'), epcs_flash_controller_0_epcs_control_port_unreg_firsttransfer, epcs_flash_controller_0_epcs_control_port_reg_firsttransfer);
  --epcs_flash_controller_0_epcs_control_port_unreg_firsttransfer first transaction, which is an e_assign
  epcs_flash_controller_0_epcs_control_port_unreg_firsttransfer <= NOT ((epcs_flash_controller_0_epcs_control_port_slavearbiterlockenable AND epcs_flash_controller_0_epcs_control_port_any_continuerequest));
  --epcs_flash_controller_0_epcs_control_port_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      epcs_flash_controller_0_epcs_control_port_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(epcs_flash_controller_0_epcs_control_port_begins_xfer) = '1' then 
        epcs_flash_controller_0_epcs_control_port_reg_firsttransfer <= epcs_flash_controller_0_epcs_control_port_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --epcs_flash_controller_0_epcs_control_port_beginbursttransfer_internal begin burst transfer, which is an e_assign
  epcs_flash_controller_0_epcs_control_port_beginbursttransfer_internal <= epcs_flash_controller_0_epcs_control_port_begins_xfer;
  --epcs_flash_controller_0_epcs_control_port_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  epcs_flash_controller_0_epcs_control_port_arbitration_holdoff_internal <= epcs_flash_controller_0_epcs_control_port_begins_xfer AND epcs_flash_controller_0_epcs_control_port_firsttransfer;
  --~epcs_flash_controller_0_epcs_control_port_read_n assignment, which is an e_mux
  epcs_flash_controller_0_epcs_control_port_read_n <= NOT ((((internal_pcp_cpu_data_master_granted_epcs_flash_controller_0_epcs_control_port AND pcp_cpu_data_master_read)) OR ((internal_pcp_cpu_instruction_master_granted_epcs_flash_controller_0_epcs_control_port AND pcp_cpu_instruction_master_read))));
  --~epcs_flash_controller_0_epcs_control_port_write_n assignment, which is an e_mux
  epcs_flash_controller_0_epcs_control_port_write_n <= NOT ((internal_pcp_cpu_data_master_granted_epcs_flash_controller_0_epcs_control_port AND pcp_cpu_data_master_write));
  shifted_address_to_epcs_flash_controller_0_epcs_control_port_from_pcp_cpu_data_master <= pcp_cpu_data_master_address_to_slave;
  --epcs_flash_controller_0_epcs_control_port_address mux, which is an e_mux
  epcs_flash_controller_0_epcs_control_port_address <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_pcp_cpu_data_master_granted_epcs_flash_controller_0_epcs_control_port)) = '1'), (A_SRL(shifted_address_to_epcs_flash_controller_0_epcs_control_port_from_pcp_cpu_data_master,std_logic_vector'("00000000000000000000000000000010"))), (A_SRL(shifted_address_to_epcs_flash_controller_0_epcs_control_port_from_pcp_cpu_instruction_master,std_logic_vector'("00000000000000000000000000000010")))), 9);
  shifted_address_to_epcs_flash_controller_0_epcs_control_port_from_pcp_cpu_instruction_master <= pcp_cpu_instruction_master_address_to_slave;
  --d1_epcs_flash_controller_0_epcs_control_port_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_epcs_flash_controller_0_epcs_control_port_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_epcs_flash_controller_0_epcs_control_port_end_xfer <= epcs_flash_controller_0_epcs_control_port_end_xfer;
    end if;

  end process;

  --epcs_flash_controller_0_epcs_control_port_waits_for_read in a cycle, which is an e_mux
  epcs_flash_controller_0_epcs_control_port_waits_for_read <= epcs_flash_controller_0_epcs_control_port_in_a_read_cycle AND epcs_flash_controller_0_epcs_control_port_begins_xfer;
  --epcs_flash_controller_0_epcs_control_port_in_a_read_cycle assignment, which is an e_assign
  epcs_flash_controller_0_epcs_control_port_in_a_read_cycle <= ((internal_pcp_cpu_data_master_granted_epcs_flash_controller_0_epcs_control_port AND pcp_cpu_data_master_read)) OR ((internal_pcp_cpu_instruction_master_granted_epcs_flash_controller_0_epcs_control_port AND pcp_cpu_instruction_master_read));
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= epcs_flash_controller_0_epcs_control_port_in_a_read_cycle;
  --epcs_flash_controller_0_epcs_control_port_waits_for_write in a cycle, which is an e_mux
  epcs_flash_controller_0_epcs_control_port_waits_for_write <= epcs_flash_controller_0_epcs_control_port_in_a_write_cycle AND epcs_flash_controller_0_epcs_control_port_begins_xfer;
  --epcs_flash_controller_0_epcs_control_port_in_a_write_cycle assignment, which is an e_assign
  epcs_flash_controller_0_epcs_control_port_in_a_write_cycle <= internal_pcp_cpu_data_master_granted_epcs_flash_controller_0_epcs_control_port AND pcp_cpu_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= epcs_flash_controller_0_epcs_control_port_in_a_write_cycle;
  wait_for_epcs_flash_controller_0_epcs_control_port_counter <= std_logic'('0');
  --assign epcs_flash_controller_0_epcs_control_port_irq_from_sa = epcs_flash_controller_0_epcs_control_port_irq so that symbol knows where to group signals which may go to master only, which is an e_assign
  epcs_flash_controller_0_epcs_control_port_irq_from_sa <= epcs_flash_controller_0_epcs_control_port_irq;
  --vhdl renameroo for output signals
  pcp_cpu_data_master_granted_epcs_flash_controller_0_epcs_control_port <= internal_pcp_cpu_data_master_granted_epcs_flash_controller_0_epcs_control_port;
  --vhdl renameroo for output signals
  pcp_cpu_data_master_qualified_request_epcs_flash_controller_0_epcs_control_port <= internal_pcp_cpu_data_master_qualified_request_epcs_flash_controller_0_epcs_control_port;
  --vhdl renameroo for output signals
  pcp_cpu_data_master_requests_epcs_flash_controller_0_epcs_control_port <= internal_pcp_cpu_data_master_requests_epcs_flash_controller_0_epcs_control_port;
  --vhdl renameroo for output signals
  pcp_cpu_instruction_master_granted_epcs_flash_controller_0_epcs_control_port <= internal_pcp_cpu_instruction_master_granted_epcs_flash_controller_0_epcs_control_port;
  --vhdl renameroo for output signals
  pcp_cpu_instruction_master_qualified_request_epcs_flash_controller_0_epcs_control_port <= internal_pcp_cpu_instruction_master_qualified_request_epcs_flash_controller_0_epcs_control_port;
  --vhdl renameroo for output signals
  pcp_cpu_instruction_master_requests_epcs_flash_controller_0_epcs_control_port <= internal_pcp_cpu_instruction_master_requests_epcs_flash_controller_0_epcs_control_port;
--synthesis translate_off
    --epcs_flash_controller_0/epcs_control_port enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --grant signals are active simultaneously, which is an e_process
    process (clk)
    VARIABLE write_line14 : line;
    begin
      if clk'event and clk = '1' then
        if (std_logic_vector'("000000000000000000000000000000") & (((std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(internal_pcp_cpu_data_master_granted_epcs_flash_controller_0_epcs_control_port))) + (std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(internal_pcp_cpu_instruction_master_granted_epcs_flash_controller_0_epcs_control_port))))))>std_logic_vector'("00000000000000000000000000000001") then 
          write(write_line14, now);
          write(write_line14, string'(": "));
          write(write_line14, string'("> 1 of grant signals are active simultaneously"));
          write(output, write_line14.all);
          deallocate (write_line14);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --saved_grant signals are active simultaneously, which is an e_process
    process (clk)
    VARIABLE write_line15 : line;
    begin
      if clk'event and clk = '1' then
        if (std_logic_vector'("000000000000000000000000000000") & (((std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(pcp_cpu_data_master_saved_grant_epcs_flash_controller_0_epcs_control_port))) + (std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(pcp_cpu_instruction_master_saved_grant_epcs_flash_controller_0_epcs_control_port))))))>std_logic_vector'("00000000000000000000000000000001") then 
          write(write_line15, now);
          write(write_line15, string'(": "));
          write(write_line15, string'("> 1 of saved_grant signals are active simultaneously"));
          write(output, write_line15.all);
          deallocate (write_line15);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity irq_gen_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal clock_crossing_0_m1_address_to_slave : IN STD_LOGIC_VECTOR (6 DOWNTO 0);
                 signal clock_crossing_0_m1_latency_counter : IN STD_LOGIC;
                 signal clock_crossing_0_m1_nativeaddress : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
                 signal clock_crossing_0_m1_read : IN STD_LOGIC;
                 signal clock_crossing_0_m1_write : IN STD_LOGIC;
                 signal clock_crossing_0_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal irq_gen_s1_readdata : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal clock_crossing_0_m1_granted_irq_gen_s1 : OUT STD_LOGIC;
                 signal clock_crossing_0_m1_qualified_request_irq_gen_s1 : OUT STD_LOGIC;
                 signal clock_crossing_0_m1_read_data_valid_irq_gen_s1 : OUT STD_LOGIC;
                 signal clock_crossing_0_m1_requests_irq_gen_s1 : OUT STD_LOGIC;
                 signal d1_irq_gen_s1_end_xfer : OUT STD_LOGIC;
                 signal irq_gen_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal irq_gen_s1_chipselect : OUT STD_LOGIC;
                 signal irq_gen_s1_readdata_from_sa : OUT STD_LOGIC;
                 signal irq_gen_s1_reset_n : OUT STD_LOGIC;
                 signal irq_gen_s1_write_n : OUT STD_LOGIC;
                 signal irq_gen_s1_writedata : OUT STD_LOGIC
              );
end entity irq_gen_s1_arbitrator;


architecture europa of irq_gen_s1_arbitrator is
                signal clock_crossing_0_m1_arbiterlock :  STD_LOGIC;
                signal clock_crossing_0_m1_arbiterlock2 :  STD_LOGIC;
                signal clock_crossing_0_m1_continuerequest :  STD_LOGIC;
                signal clock_crossing_0_m1_saved_grant_irq_gen_s1 :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_irq_gen_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_clock_crossing_0_m1_granted_irq_gen_s1 :  STD_LOGIC;
                signal internal_clock_crossing_0_m1_qualified_request_irq_gen_s1 :  STD_LOGIC;
                signal internal_clock_crossing_0_m1_requests_irq_gen_s1 :  STD_LOGIC;
                signal irq_gen_s1_allgrants :  STD_LOGIC;
                signal irq_gen_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal irq_gen_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal irq_gen_s1_any_continuerequest :  STD_LOGIC;
                signal irq_gen_s1_arb_counter_enable :  STD_LOGIC;
                signal irq_gen_s1_arb_share_counter :  STD_LOGIC;
                signal irq_gen_s1_arb_share_counter_next_value :  STD_LOGIC;
                signal irq_gen_s1_arb_share_set_values :  STD_LOGIC;
                signal irq_gen_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal irq_gen_s1_begins_xfer :  STD_LOGIC;
                signal irq_gen_s1_end_xfer :  STD_LOGIC;
                signal irq_gen_s1_firsttransfer :  STD_LOGIC;
                signal irq_gen_s1_grant_vector :  STD_LOGIC;
                signal irq_gen_s1_in_a_read_cycle :  STD_LOGIC;
                signal irq_gen_s1_in_a_write_cycle :  STD_LOGIC;
                signal irq_gen_s1_master_qreq_vector :  STD_LOGIC;
                signal irq_gen_s1_non_bursting_master_requests :  STD_LOGIC;
                signal irq_gen_s1_reg_firsttransfer :  STD_LOGIC;
                signal irq_gen_s1_slavearbiterlockenable :  STD_LOGIC;
                signal irq_gen_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal irq_gen_s1_unreg_firsttransfer :  STD_LOGIC;
                signal irq_gen_s1_waits_for_read :  STD_LOGIC;
                signal irq_gen_s1_waits_for_write :  STD_LOGIC;
                signal wait_for_irq_gen_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT irq_gen_s1_end_xfer;
    end if;

  end process;

  irq_gen_s1_begins_xfer <= NOT d1_reasons_to_wait AND (internal_clock_crossing_0_m1_qualified_request_irq_gen_s1);
  --assign irq_gen_s1_readdata_from_sa = irq_gen_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  irq_gen_s1_readdata_from_sa <= irq_gen_s1_readdata;
  internal_clock_crossing_0_m1_requests_irq_gen_s1 <= to_std_logic(((Std_Logic_Vector'(clock_crossing_0_m1_address_to_slave(6 DOWNTO 4) & std_logic_vector'("0000")) = std_logic_vector'("1000000")))) AND ((clock_crossing_0_m1_read OR clock_crossing_0_m1_write));
  --irq_gen_s1_arb_share_counter set values, which is an e_mux
  irq_gen_s1_arb_share_set_values <= std_logic'('1');
  --irq_gen_s1_non_bursting_master_requests mux, which is an e_mux
  irq_gen_s1_non_bursting_master_requests <= internal_clock_crossing_0_m1_requests_irq_gen_s1;
  --irq_gen_s1_any_bursting_master_saved_grant mux, which is an e_mux
  irq_gen_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --irq_gen_s1_arb_share_counter_next_value assignment, which is an e_assign
  irq_gen_s1_arb_share_counter_next_value <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(irq_gen_s1_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(irq_gen_s1_arb_share_set_values))) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(irq_gen_s1_arb_share_counter) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(irq_gen_s1_arb_share_counter))) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))));
  --irq_gen_s1_allgrants all slave grants, which is an e_mux
  irq_gen_s1_allgrants <= irq_gen_s1_grant_vector;
  --irq_gen_s1_end_xfer assignment, which is an e_assign
  irq_gen_s1_end_xfer <= NOT ((irq_gen_s1_waits_for_read OR irq_gen_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_irq_gen_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_irq_gen_s1 <= irq_gen_s1_end_xfer AND (((NOT irq_gen_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --irq_gen_s1_arb_share_counter arbitration counter enable, which is an e_assign
  irq_gen_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_irq_gen_s1 AND irq_gen_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_irq_gen_s1 AND NOT irq_gen_s1_non_bursting_master_requests));
  --irq_gen_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      irq_gen_s1_arb_share_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(irq_gen_s1_arb_counter_enable) = '1' then 
        irq_gen_s1_arb_share_counter <= irq_gen_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --irq_gen_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      irq_gen_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((irq_gen_s1_master_qreq_vector AND end_xfer_arb_share_counter_term_irq_gen_s1)) OR ((end_xfer_arb_share_counter_term_irq_gen_s1 AND NOT irq_gen_s1_non_bursting_master_requests)))) = '1' then 
        irq_gen_s1_slavearbiterlockenable <= irq_gen_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --clock_crossing_0/m1 irq_gen/s1 arbiterlock, which is an e_assign
  clock_crossing_0_m1_arbiterlock <= irq_gen_s1_slavearbiterlockenable AND clock_crossing_0_m1_continuerequest;
  --irq_gen_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  irq_gen_s1_slavearbiterlockenable2 <= irq_gen_s1_arb_share_counter_next_value;
  --clock_crossing_0/m1 irq_gen/s1 arbiterlock2, which is an e_assign
  clock_crossing_0_m1_arbiterlock2 <= irq_gen_s1_slavearbiterlockenable2 AND clock_crossing_0_m1_continuerequest;
  --irq_gen_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  irq_gen_s1_any_continuerequest <= std_logic'('1');
  --clock_crossing_0_m1_continuerequest continued request, which is an e_assign
  clock_crossing_0_m1_continuerequest <= std_logic'('1');
  internal_clock_crossing_0_m1_qualified_request_irq_gen_s1 <= internal_clock_crossing_0_m1_requests_irq_gen_s1 AND NOT ((clock_crossing_0_m1_read AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(clock_crossing_0_m1_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))))));
  --local readdatavalid clock_crossing_0_m1_read_data_valid_irq_gen_s1, which is an e_mux
  clock_crossing_0_m1_read_data_valid_irq_gen_s1 <= (internal_clock_crossing_0_m1_granted_irq_gen_s1 AND clock_crossing_0_m1_read) AND NOT irq_gen_s1_waits_for_read;
  --irq_gen_s1_writedata mux, which is an e_mux
  irq_gen_s1_writedata <= clock_crossing_0_m1_writedata(0);
  --master is always granted when requested
  internal_clock_crossing_0_m1_granted_irq_gen_s1 <= internal_clock_crossing_0_m1_qualified_request_irq_gen_s1;
  --clock_crossing_0/m1 saved-grant irq_gen/s1, which is an e_assign
  clock_crossing_0_m1_saved_grant_irq_gen_s1 <= internal_clock_crossing_0_m1_requests_irq_gen_s1;
  --allow new arb cycle for irq_gen/s1, which is an e_assign
  irq_gen_s1_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  irq_gen_s1_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  irq_gen_s1_master_qreq_vector <= std_logic'('1');
  --irq_gen_s1_reset_n assignment, which is an e_assign
  irq_gen_s1_reset_n <= reset_n;
  irq_gen_s1_chipselect <= internal_clock_crossing_0_m1_granted_irq_gen_s1;
  --irq_gen_s1_firsttransfer first transaction, which is an e_assign
  irq_gen_s1_firsttransfer <= A_WE_StdLogic((std_logic'(irq_gen_s1_begins_xfer) = '1'), irq_gen_s1_unreg_firsttransfer, irq_gen_s1_reg_firsttransfer);
  --irq_gen_s1_unreg_firsttransfer first transaction, which is an e_assign
  irq_gen_s1_unreg_firsttransfer <= NOT ((irq_gen_s1_slavearbiterlockenable AND irq_gen_s1_any_continuerequest));
  --irq_gen_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      irq_gen_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(irq_gen_s1_begins_xfer) = '1' then 
        irq_gen_s1_reg_firsttransfer <= irq_gen_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --irq_gen_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  irq_gen_s1_beginbursttransfer_internal <= irq_gen_s1_begins_xfer;
  --~irq_gen_s1_write_n assignment, which is an e_mux
  irq_gen_s1_write_n <= NOT ((internal_clock_crossing_0_m1_granted_irq_gen_s1 AND clock_crossing_0_m1_write));
  --irq_gen_s1_address mux, which is an e_mux
  irq_gen_s1_address <= clock_crossing_0_m1_nativeaddress (1 DOWNTO 0);
  --d1_irq_gen_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_irq_gen_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_irq_gen_s1_end_xfer <= irq_gen_s1_end_xfer;
    end if;

  end process;

  --irq_gen_s1_waits_for_read in a cycle, which is an e_mux
  irq_gen_s1_waits_for_read <= irq_gen_s1_in_a_read_cycle AND irq_gen_s1_begins_xfer;
  --irq_gen_s1_in_a_read_cycle assignment, which is an e_assign
  irq_gen_s1_in_a_read_cycle <= internal_clock_crossing_0_m1_granted_irq_gen_s1 AND clock_crossing_0_m1_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= irq_gen_s1_in_a_read_cycle;
  --irq_gen_s1_waits_for_write in a cycle, which is an e_mux
  irq_gen_s1_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(irq_gen_s1_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --irq_gen_s1_in_a_write_cycle assignment, which is an e_assign
  irq_gen_s1_in_a_write_cycle <= internal_clock_crossing_0_m1_granted_irq_gen_s1 AND clock_crossing_0_m1_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= irq_gen_s1_in_a_write_cycle;
  wait_for_irq_gen_s1_counter <= std_logic'('0');
  --vhdl renameroo for output signals
  clock_crossing_0_m1_granted_irq_gen_s1 <= internal_clock_crossing_0_m1_granted_irq_gen_s1;
  --vhdl renameroo for output signals
  clock_crossing_0_m1_qualified_request_irq_gen_s1 <= internal_clock_crossing_0_m1_qualified_request_irq_gen_s1;
  --vhdl renameroo for output signals
  clock_crossing_0_m1_requests_irq_gen_s1 <= internal_clock_crossing_0_m1_requests_irq_gen_s1;
--synthesis translate_off
    --irq_gen/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity jtag_uart_0_avalon_jtag_slave_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal jtag_uart_0_avalon_jtag_slave_dataavailable : IN STD_LOGIC;
                 signal jtag_uart_0_avalon_jtag_slave_irq : IN STD_LOGIC;
                 signal jtag_uart_0_avalon_jtag_slave_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal jtag_uart_0_avalon_jtag_slave_readyfordata : IN STD_LOGIC;
                 signal jtag_uart_0_avalon_jtag_slave_waitrequest : IN STD_LOGIC;
                 signal niosII_openMac_clock_0_out_address_to_slave : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal niosII_openMac_clock_0_out_nativeaddress : IN STD_LOGIC;
                 signal niosII_openMac_clock_0_out_read : IN STD_LOGIC;
                 signal niosII_openMac_clock_0_out_write : IN STD_LOGIC;
                 signal niosII_openMac_clock_0_out_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal d1_jtag_uart_0_avalon_jtag_slave_end_xfer : OUT STD_LOGIC;
                 signal jtag_uart_0_avalon_jtag_slave_address : OUT STD_LOGIC;
                 signal jtag_uart_0_avalon_jtag_slave_chipselect : OUT STD_LOGIC;
                 signal jtag_uart_0_avalon_jtag_slave_dataavailable_from_sa : OUT STD_LOGIC;
                 signal jtag_uart_0_avalon_jtag_slave_irq_from_sa : OUT STD_LOGIC;
                 signal jtag_uart_0_avalon_jtag_slave_read_n : OUT STD_LOGIC;
                 signal jtag_uart_0_avalon_jtag_slave_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal jtag_uart_0_avalon_jtag_slave_readyfordata_from_sa : OUT STD_LOGIC;
                 signal jtag_uart_0_avalon_jtag_slave_reset_n : OUT STD_LOGIC;
                 signal jtag_uart_0_avalon_jtag_slave_waitrequest_from_sa : OUT STD_LOGIC;
                 signal jtag_uart_0_avalon_jtag_slave_write_n : OUT STD_LOGIC;
                 signal jtag_uart_0_avalon_jtag_slave_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal niosII_openMac_clock_0_out_granted_jtag_uart_0_avalon_jtag_slave : OUT STD_LOGIC;
                 signal niosII_openMac_clock_0_out_qualified_request_jtag_uart_0_avalon_jtag_slave : OUT STD_LOGIC;
                 signal niosII_openMac_clock_0_out_read_data_valid_jtag_uart_0_avalon_jtag_slave : OUT STD_LOGIC;
                 signal niosII_openMac_clock_0_out_requests_jtag_uart_0_avalon_jtag_slave : OUT STD_LOGIC
              );
end entity jtag_uart_0_avalon_jtag_slave_arbitrator;


architecture europa of jtag_uart_0_avalon_jtag_slave_arbitrator is
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_jtag_uart_0_avalon_jtag_slave :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_jtag_uart_0_avalon_jtag_slave_waitrequest_from_sa :  STD_LOGIC;
                signal internal_niosII_openMac_clock_0_out_granted_jtag_uart_0_avalon_jtag_slave :  STD_LOGIC;
                signal internal_niosII_openMac_clock_0_out_qualified_request_jtag_uart_0_avalon_jtag_slave :  STD_LOGIC;
                signal internal_niosII_openMac_clock_0_out_requests_jtag_uart_0_avalon_jtag_slave :  STD_LOGIC;
                signal jtag_uart_0_avalon_jtag_slave_allgrants :  STD_LOGIC;
                signal jtag_uart_0_avalon_jtag_slave_allow_new_arb_cycle :  STD_LOGIC;
                signal jtag_uart_0_avalon_jtag_slave_any_bursting_master_saved_grant :  STD_LOGIC;
                signal jtag_uart_0_avalon_jtag_slave_any_continuerequest :  STD_LOGIC;
                signal jtag_uart_0_avalon_jtag_slave_arb_counter_enable :  STD_LOGIC;
                signal jtag_uart_0_avalon_jtag_slave_arb_share_counter :  STD_LOGIC;
                signal jtag_uart_0_avalon_jtag_slave_arb_share_counter_next_value :  STD_LOGIC;
                signal jtag_uart_0_avalon_jtag_slave_arb_share_set_values :  STD_LOGIC;
                signal jtag_uart_0_avalon_jtag_slave_beginbursttransfer_internal :  STD_LOGIC;
                signal jtag_uart_0_avalon_jtag_slave_begins_xfer :  STD_LOGIC;
                signal jtag_uart_0_avalon_jtag_slave_end_xfer :  STD_LOGIC;
                signal jtag_uart_0_avalon_jtag_slave_firsttransfer :  STD_LOGIC;
                signal jtag_uart_0_avalon_jtag_slave_grant_vector :  STD_LOGIC;
                signal jtag_uart_0_avalon_jtag_slave_in_a_read_cycle :  STD_LOGIC;
                signal jtag_uart_0_avalon_jtag_slave_in_a_write_cycle :  STD_LOGIC;
                signal jtag_uart_0_avalon_jtag_slave_master_qreq_vector :  STD_LOGIC;
                signal jtag_uart_0_avalon_jtag_slave_non_bursting_master_requests :  STD_LOGIC;
                signal jtag_uart_0_avalon_jtag_slave_reg_firsttransfer :  STD_LOGIC;
                signal jtag_uart_0_avalon_jtag_slave_slavearbiterlockenable :  STD_LOGIC;
                signal jtag_uart_0_avalon_jtag_slave_slavearbiterlockenable2 :  STD_LOGIC;
                signal jtag_uart_0_avalon_jtag_slave_unreg_firsttransfer :  STD_LOGIC;
                signal jtag_uart_0_avalon_jtag_slave_waits_for_read :  STD_LOGIC;
                signal jtag_uart_0_avalon_jtag_slave_waits_for_write :  STD_LOGIC;
                signal niosII_openMac_clock_0_out_arbiterlock :  STD_LOGIC;
                signal niosII_openMac_clock_0_out_arbiterlock2 :  STD_LOGIC;
                signal niosII_openMac_clock_0_out_continuerequest :  STD_LOGIC;
                signal niosII_openMac_clock_0_out_saved_grant_jtag_uart_0_avalon_jtag_slave :  STD_LOGIC;
                signal wait_for_jtag_uart_0_avalon_jtag_slave_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT jtag_uart_0_avalon_jtag_slave_end_xfer;
    end if;

  end process;

  jtag_uart_0_avalon_jtag_slave_begins_xfer <= NOT d1_reasons_to_wait AND (internal_niosII_openMac_clock_0_out_qualified_request_jtag_uart_0_avalon_jtag_slave);
  --assign jtag_uart_0_avalon_jtag_slave_readdata_from_sa = jtag_uart_0_avalon_jtag_slave_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  jtag_uart_0_avalon_jtag_slave_readdata_from_sa <= jtag_uart_0_avalon_jtag_slave_readdata;
  internal_niosII_openMac_clock_0_out_requests_jtag_uart_0_avalon_jtag_slave <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((niosII_openMac_clock_0_out_read OR niosII_openMac_clock_0_out_write)))))));
  --assign jtag_uart_0_avalon_jtag_slave_dataavailable_from_sa = jtag_uart_0_avalon_jtag_slave_dataavailable so that symbol knows where to group signals which may go to master only, which is an e_assign
  jtag_uart_0_avalon_jtag_slave_dataavailable_from_sa <= jtag_uart_0_avalon_jtag_slave_dataavailable;
  --assign jtag_uart_0_avalon_jtag_slave_readyfordata_from_sa = jtag_uart_0_avalon_jtag_slave_readyfordata so that symbol knows where to group signals which may go to master only, which is an e_assign
  jtag_uart_0_avalon_jtag_slave_readyfordata_from_sa <= jtag_uart_0_avalon_jtag_slave_readyfordata;
  --assign jtag_uart_0_avalon_jtag_slave_waitrequest_from_sa = jtag_uart_0_avalon_jtag_slave_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_jtag_uart_0_avalon_jtag_slave_waitrequest_from_sa <= jtag_uart_0_avalon_jtag_slave_waitrequest;
  --jtag_uart_0_avalon_jtag_slave_arb_share_counter set values, which is an e_mux
  jtag_uart_0_avalon_jtag_slave_arb_share_set_values <= std_logic'('1');
  --jtag_uart_0_avalon_jtag_slave_non_bursting_master_requests mux, which is an e_mux
  jtag_uart_0_avalon_jtag_slave_non_bursting_master_requests <= internal_niosII_openMac_clock_0_out_requests_jtag_uart_0_avalon_jtag_slave;
  --jtag_uart_0_avalon_jtag_slave_any_bursting_master_saved_grant mux, which is an e_mux
  jtag_uart_0_avalon_jtag_slave_any_bursting_master_saved_grant <= std_logic'('0');
  --jtag_uart_0_avalon_jtag_slave_arb_share_counter_next_value assignment, which is an e_assign
  jtag_uart_0_avalon_jtag_slave_arb_share_counter_next_value <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(jtag_uart_0_avalon_jtag_slave_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(jtag_uart_0_avalon_jtag_slave_arb_share_set_values))) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(jtag_uart_0_avalon_jtag_slave_arb_share_counter) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(jtag_uart_0_avalon_jtag_slave_arb_share_counter))) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))));
  --jtag_uart_0_avalon_jtag_slave_allgrants all slave grants, which is an e_mux
  jtag_uart_0_avalon_jtag_slave_allgrants <= jtag_uart_0_avalon_jtag_slave_grant_vector;
  --jtag_uart_0_avalon_jtag_slave_end_xfer assignment, which is an e_assign
  jtag_uart_0_avalon_jtag_slave_end_xfer <= NOT ((jtag_uart_0_avalon_jtag_slave_waits_for_read OR jtag_uart_0_avalon_jtag_slave_waits_for_write));
  --end_xfer_arb_share_counter_term_jtag_uart_0_avalon_jtag_slave arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_jtag_uart_0_avalon_jtag_slave <= jtag_uart_0_avalon_jtag_slave_end_xfer AND (((NOT jtag_uart_0_avalon_jtag_slave_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --jtag_uart_0_avalon_jtag_slave_arb_share_counter arbitration counter enable, which is an e_assign
  jtag_uart_0_avalon_jtag_slave_arb_counter_enable <= ((end_xfer_arb_share_counter_term_jtag_uart_0_avalon_jtag_slave AND jtag_uart_0_avalon_jtag_slave_allgrants)) OR ((end_xfer_arb_share_counter_term_jtag_uart_0_avalon_jtag_slave AND NOT jtag_uart_0_avalon_jtag_slave_non_bursting_master_requests));
  --jtag_uart_0_avalon_jtag_slave_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      jtag_uart_0_avalon_jtag_slave_arb_share_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(jtag_uart_0_avalon_jtag_slave_arb_counter_enable) = '1' then 
        jtag_uart_0_avalon_jtag_slave_arb_share_counter <= jtag_uart_0_avalon_jtag_slave_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --jtag_uart_0_avalon_jtag_slave_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      jtag_uart_0_avalon_jtag_slave_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((jtag_uart_0_avalon_jtag_slave_master_qreq_vector AND end_xfer_arb_share_counter_term_jtag_uart_0_avalon_jtag_slave)) OR ((end_xfer_arb_share_counter_term_jtag_uart_0_avalon_jtag_slave AND NOT jtag_uart_0_avalon_jtag_slave_non_bursting_master_requests)))) = '1' then 
        jtag_uart_0_avalon_jtag_slave_slavearbiterlockenable <= jtag_uart_0_avalon_jtag_slave_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --niosII_openMac_clock_0/out jtag_uart_0/avalon_jtag_slave arbiterlock, which is an e_assign
  niosII_openMac_clock_0_out_arbiterlock <= jtag_uart_0_avalon_jtag_slave_slavearbiterlockenable AND niosII_openMac_clock_0_out_continuerequest;
  --jtag_uart_0_avalon_jtag_slave_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  jtag_uart_0_avalon_jtag_slave_slavearbiterlockenable2 <= jtag_uart_0_avalon_jtag_slave_arb_share_counter_next_value;
  --niosII_openMac_clock_0/out jtag_uart_0/avalon_jtag_slave arbiterlock2, which is an e_assign
  niosII_openMac_clock_0_out_arbiterlock2 <= jtag_uart_0_avalon_jtag_slave_slavearbiterlockenable2 AND niosII_openMac_clock_0_out_continuerequest;
  --jtag_uart_0_avalon_jtag_slave_any_continuerequest at least one master continues requesting, which is an e_assign
  jtag_uart_0_avalon_jtag_slave_any_continuerequest <= std_logic'('1');
  --niosII_openMac_clock_0_out_continuerequest continued request, which is an e_assign
  niosII_openMac_clock_0_out_continuerequest <= std_logic'('1');
  internal_niosII_openMac_clock_0_out_qualified_request_jtag_uart_0_avalon_jtag_slave <= internal_niosII_openMac_clock_0_out_requests_jtag_uart_0_avalon_jtag_slave;
  --jtag_uart_0_avalon_jtag_slave_writedata mux, which is an e_mux
  jtag_uart_0_avalon_jtag_slave_writedata <= niosII_openMac_clock_0_out_writedata;
  --master is always granted when requested
  internal_niosII_openMac_clock_0_out_granted_jtag_uart_0_avalon_jtag_slave <= internal_niosII_openMac_clock_0_out_qualified_request_jtag_uart_0_avalon_jtag_slave;
  --niosII_openMac_clock_0/out saved-grant jtag_uart_0/avalon_jtag_slave, which is an e_assign
  niosII_openMac_clock_0_out_saved_grant_jtag_uart_0_avalon_jtag_slave <= internal_niosII_openMac_clock_0_out_requests_jtag_uart_0_avalon_jtag_slave;
  --allow new arb cycle for jtag_uart_0/avalon_jtag_slave, which is an e_assign
  jtag_uart_0_avalon_jtag_slave_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  jtag_uart_0_avalon_jtag_slave_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  jtag_uart_0_avalon_jtag_slave_master_qreq_vector <= std_logic'('1');
  --jtag_uart_0_avalon_jtag_slave_reset_n assignment, which is an e_assign
  jtag_uart_0_avalon_jtag_slave_reset_n <= reset_n;
  jtag_uart_0_avalon_jtag_slave_chipselect <= internal_niosII_openMac_clock_0_out_granted_jtag_uart_0_avalon_jtag_slave;
  --jtag_uart_0_avalon_jtag_slave_firsttransfer first transaction, which is an e_assign
  jtag_uart_0_avalon_jtag_slave_firsttransfer <= A_WE_StdLogic((std_logic'(jtag_uart_0_avalon_jtag_slave_begins_xfer) = '1'), jtag_uart_0_avalon_jtag_slave_unreg_firsttransfer, jtag_uart_0_avalon_jtag_slave_reg_firsttransfer);
  --jtag_uart_0_avalon_jtag_slave_unreg_firsttransfer first transaction, which is an e_assign
  jtag_uart_0_avalon_jtag_slave_unreg_firsttransfer <= NOT ((jtag_uart_0_avalon_jtag_slave_slavearbiterlockenable AND jtag_uart_0_avalon_jtag_slave_any_continuerequest));
  --jtag_uart_0_avalon_jtag_slave_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      jtag_uart_0_avalon_jtag_slave_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(jtag_uart_0_avalon_jtag_slave_begins_xfer) = '1' then 
        jtag_uart_0_avalon_jtag_slave_reg_firsttransfer <= jtag_uart_0_avalon_jtag_slave_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --jtag_uart_0_avalon_jtag_slave_beginbursttransfer_internal begin burst transfer, which is an e_assign
  jtag_uart_0_avalon_jtag_slave_beginbursttransfer_internal <= jtag_uart_0_avalon_jtag_slave_begins_xfer;
  --~jtag_uart_0_avalon_jtag_slave_read_n assignment, which is an e_mux
  jtag_uart_0_avalon_jtag_slave_read_n <= NOT ((internal_niosII_openMac_clock_0_out_granted_jtag_uart_0_avalon_jtag_slave AND niosII_openMac_clock_0_out_read));
  --~jtag_uart_0_avalon_jtag_slave_write_n assignment, which is an e_mux
  jtag_uart_0_avalon_jtag_slave_write_n <= NOT ((internal_niosII_openMac_clock_0_out_granted_jtag_uart_0_avalon_jtag_slave AND niosII_openMac_clock_0_out_write));
  --jtag_uart_0_avalon_jtag_slave_address mux, which is an e_mux
  jtag_uart_0_avalon_jtag_slave_address <= niosII_openMac_clock_0_out_nativeaddress;
  --d1_jtag_uart_0_avalon_jtag_slave_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_jtag_uart_0_avalon_jtag_slave_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_jtag_uart_0_avalon_jtag_slave_end_xfer <= jtag_uart_0_avalon_jtag_slave_end_xfer;
    end if;

  end process;

  --jtag_uart_0_avalon_jtag_slave_waits_for_read in a cycle, which is an e_mux
  jtag_uart_0_avalon_jtag_slave_waits_for_read <= jtag_uart_0_avalon_jtag_slave_in_a_read_cycle AND internal_jtag_uart_0_avalon_jtag_slave_waitrequest_from_sa;
  --jtag_uart_0_avalon_jtag_slave_in_a_read_cycle assignment, which is an e_assign
  jtag_uart_0_avalon_jtag_slave_in_a_read_cycle <= internal_niosII_openMac_clock_0_out_granted_jtag_uart_0_avalon_jtag_slave AND niosII_openMac_clock_0_out_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= jtag_uart_0_avalon_jtag_slave_in_a_read_cycle;
  --jtag_uart_0_avalon_jtag_slave_waits_for_write in a cycle, which is an e_mux
  jtag_uart_0_avalon_jtag_slave_waits_for_write <= jtag_uart_0_avalon_jtag_slave_in_a_write_cycle AND internal_jtag_uart_0_avalon_jtag_slave_waitrequest_from_sa;
  --jtag_uart_0_avalon_jtag_slave_in_a_write_cycle assignment, which is an e_assign
  jtag_uart_0_avalon_jtag_slave_in_a_write_cycle <= internal_niosII_openMac_clock_0_out_granted_jtag_uart_0_avalon_jtag_slave AND niosII_openMac_clock_0_out_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= jtag_uart_0_avalon_jtag_slave_in_a_write_cycle;
  wait_for_jtag_uart_0_avalon_jtag_slave_counter <= std_logic'('0');
  --assign jtag_uart_0_avalon_jtag_slave_irq_from_sa = jtag_uart_0_avalon_jtag_slave_irq so that symbol knows where to group signals which may go to master only, which is an e_assign
  jtag_uart_0_avalon_jtag_slave_irq_from_sa <= jtag_uart_0_avalon_jtag_slave_irq;
  --vhdl renameroo for output signals
  jtag_uart_0_avalon_jtag_slave_waitrequest_from_sa <= internal_jtag_uart_0_avalon_jtag_slave_waitrequest_from_sa;
  --vhdl renameroo for output signals
  niosII_openMac_clock_0_out_granted_jtag_uart_0_avalon_jtag_slave <= internal_niosII_openMac_clock_0_out_granted_jtag_uart_0_avalon_jtag_slave;
  --vhdl renameroo for output signals
  niosII_openMac_clock_0_out_qualified_request_jtag_uart_0_avalon_jtag_slave <= internal_niosII_openMac_clock_0_out_qualified_request_jtag_uart_0_avalon_jtag_slave;
  --vhdl renameroo for output signals
  niosII_openMac_clock_0_out_requests_jtag_uart_0_avalon_jtag_slave <= internal_niosII_openMac_clock_0_out_requests_jtag_uart_0_avalon_jtag_slave;
--synthesis translate_off
    --jtag_uart_0/avalon_jtag_slave enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity jtag_uart_1_avalon_jtag_slave_arbitrator is 
        port (
              -- inputs:
                 signal ap_cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (25 DOWNTO 0);
                 signal ap_cpu_data_master_read : IN STD_LOGIC;
                 signal ap_cpu_data_master_waitrequest : IN STD_LOGIC;
                 signal ap_cpu_data_master_write : IN STD_LOGIC;
                 signal ap_cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal clk : IN STD_LOGIC;
                 signal jtag_uart_1_avalon_jtag_slave_dataavailable : IN STD_LOGIC;
                 signal jtag_uart_1_avalon_jtag_slave_irq : IN STD_LOGIC;
                 signal jtag_uart_1_avalon_jtag_slave_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal jtag_uart_1_avalon_jtag_slave_readyfordata : IN STD_LOGIC;
                 signal jtag_uart_1_avalon_jtag_slave_waitrequest : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal ap_cpu_data_master_granted_jtag_uart_1_avalon_jtag_slave : OUT STD_LOGIC;
                 signal ap_cpu_data_master_qualified_request_jtag_uart_1_avalon_jtag_slave : OUT STD_LOGIC;
                 signal ap_cpu_data_master_read_data_valid_jtag_uart_1_avalon_jtag_slave : OUT STD_LOGIC;
                 signal ap_cpu_data_master_requests_jtag_uart_1_avalon_jtag_slave : OUT STD_LOGIC;
                 signal d1_jtag_uart_1_avalon_jtag_slave_end_xfer : OUT STD_LOGIC;
                 signal jtag_uart_1_avalon_jtag_slave_address : OUT STD_LOGIC;
                 signal jtag_uart_1_avalon_jtag_slave_chipselect : OUT STD_LOGIC;
                 signal jtag_uart_1_avalon_jtag_slave_dataavailable_from_sa : OUT STD_LOGIC;
                 signal jtag_uart_1_avalon_jtag_slave_irq_from_sa : OUT STD_LOGIC;
                 signal jtag_uart_1_avalon_jtag_slave_read_n : OUT STD_LOGIC;
                 signal jtag_uart_1_avalon_jtag_slave_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal jtag_uart_1_avalon_jtag_slave_readyfordata_from_sa : OUT STD_LOGIC;
                 signal jtag_uart_1_avalon_jtag_slave_reset_n : OUT STD_LOGIC;
                 signal jtag_uart_1_avalon_jtag_slave_waitrequest_from_sa : OUT STD_LOGIC;
                 signal jtag_uart_1_avalon_jtag_slave_write_n : OUT STD_LOGIC;
                 signal jtag_uart_1_avalon_jtag_slave_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
              );
end entity jtag_uart_1_avalon_jtag_slave_arbitrator;


architecture europa of jtag_uart_1_avalon_jtag_slave_arbitrator is
                signal ap_cpu_data_master_arbiterlock :  STD_LOGIC;
                signal ap_cpu_data_master_arbiterlock2 :  STD_LOGIC;
                signal ap_cpu_data_master_continuerequest :  STD_LOGIC;
                signal ap_cpu_data_master_saved_grant_jtag_uart_1_avalon_jtag_slave :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_jtag_uart_1_avalon_jtag_slave :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_ap_cpu_data_master_granted_jtag_uart_1_avalon_jtag_slave :  STD_LOGIC;
                signal internal_ap_cpu_data_master_qualified_request_jtag_uart_1_avalon_jtag_slave :  STD_LOGIC;
                signal internal_ap_cpu_data_master_requests_jtag_uart_1_avalon_jtag_slave :  STD_LOGIC;
                signal internal_jtag_uart_1_avalon_jtag_slave_waitrequest_from_sa :  STD_LOGIC;
                signal jtag_uart_1_avalon_jtag_slave_allgrants :  STD_LOGIC;
                signal jtag_uart_1_avalon_jtag_slave_allow_new_arb_cycle :  STD_LOGIC;
                signal jtag_uart_1_avalon_jtag_slave_any_bursting_master_saved_grant :  STD_LOGIC;
                signal jtag_uart_1_avalon_jtag_slave_any_continuerequest :  STD_LOGIC;
                signal jtag_uart_1_avalon_jtag_slave_arb_counter_enable :  STD_LOGIC;
                signal jtag_uart_1_avalon_jtag_slave_arb_share_counter :  STD_LOGIC;
                signal jtag_uart_1_avalon_jtag_slave_arb_share_counter_next_value :  STD_LOGIC;
                signal jtag_uart_1_avalon_jtag_slave_arb_share_set_values :  STD_LOGIC;
                signal jtag_uart_1_avalon_jtag_slave_beginbursttransfer_internal :  STD_LOGIC;
                signal jtag_uart_1_avalon_jtag_slave_begins_xfer :  STD_LOGIC;
                signal jtag_uart_1_avalon_jtag_slave_end_xfer :  STD_LOGIC;
                signal jtag_uart_1_avalon_jtag_slave_firsttransfer :  STD_LOGIC;
                signal jtag_uart_1_avalon_jtag_slave_grant_vector :  STD_LOGIC;
                signal jtag_uart_1_avalon_jtag_slave_in_a_read_cycle :  STD_LOGIC;
                signal jtag_uart_1_avalon_jtag_slave_in_a_write_cycle :  STD_LOGIC;
                signal jtag_uart_1_avalon_jtag_slave_master_qreq_vector :  STD_LOGIC;
                signal jtag_uart_1_avalon_jtag_slave_non_bursting_master_requests :  STD_LOGIC;
                signal jtag_uart_1_avalon_jtag_slave_reg_firsttransfer :  STD_LOGIC;
                signal jtag_uart_1_avalon_jtag_slave_slavearbiterlockenable :  STD_LOGIC;
                signal jtag_uart_1_avalon_jtag_slave_slavearbiterlockenable2 :  STD_LOGIC;
                signal jtag_uart_1_avalon_jtag_slave_unreg_firsttransfer :  STD_LOGIC;
                signal jtag_uart_1_avalon_jtag_slave_waits_for_read :  STD_LOGIC;
                signal jtag_uart_1_avalon_jtag_slave_waits_for_write :  STD_LOGIC;
                signal shifted_address_to_jtag_uart_1_avalon_jtag_slave_from_ap_cpu_data_master :  STD_LOGIC_VECTOR (25 DOWNTO 0);
                signal wait_for_jtag_uart_1_avalon_jtag_slave_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT jtag_uart_1_avalon_jtag_slave_end_xfer;
    end if;

  end process;

  jtag_uart_1_avalon_jtag_slave_begins_xfer <= NOT d1_reasons_to_wait AND (internal_ap_cpu_data_master_qualified_request_jtag_uart_1_avalon_jtag_slave);
  --assign jtag_uart_1_avalon_jtag_slave_readdata_from_sa = jtag_uart_1_avalon_jtag_slave_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  jtag_uart_1_avalon_jtag_slave_readdata_from_sa <= jtag_uart_1_avalon_jtag_slave_readdata;
  internal_ap_cpu_data_master_requests_jtag_uart_1_avalon_jtag_slave <= to_std_logic(((Std_Logic_Vector'(ap_cpu_data_master_address_to_slave(25 DOWNTO 3) & std_logic_vector'("000")) = std_logic_vector'("11000000100001000000000000")))) AND ((ap_cpu_data_master_read OR ap_cpu_data_master_write));
  --assign jtag_uart_1_avalon_jtag_slave_dataavailable_from_sa = jtag_uart_1_avalon_jtag_slave_dataavailable so that symbol knows where to group signals which may go to master only, which is an e_assign
  jtag_uart_1_avalon_jtag_slave_dataavailable_from_sa <= jtag_uart_1_avalon_jtag_slave_dataavailable;
  --assign jtag_uart_1_avalon_jtag_slave_readyfordata_from_sa = jtag_uart_1_avalon_jtag_slave_readyfordata so that symbol knows where to group signals which may go to master only, which is an e_assign
  jtag_uart_1_avalon_jtag_slave_readyfordata_from_sa <= jtag_uart_1_avalon_jtag_slave_readyfordata;
  --assign jtag_uart_1_avalon_jtag_slave_waitrequest_from_sa = jtag_uart_1_avalon_jtag_slave_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_jtag_uart_1_avalon_jtag_slave_waitrequest_from_sa <= jtag_uart_1_avalon_jtag_slave_waitrequest;
  --jtag_uart_1_avalon_jtag_slave_arb_share_counter set values, which is an e_mux
  jtag_uart_1_avalon_jtag_slave_arb_share_set_values <= std_logic'('1');
  --jtag_uart_1_avalon_jtag_slave_non_bursting_master_requests mux, which is an e_mux
  jtag_uart_1_avalon_jtag_slave_non_bursting_master_requests <= internal_ap_cpu_data_master_requests_jtag_uart_1_avalon_jtag_slave;
  --jtag_uart_1_avalon_jtag_slave_any_bursting_master_saved_grant mux, which is an e_mux
  jtag_uart_1_avalon_jtag_slave_any_bursting_master_saved_grant <= std_logic'('0');
  --jtag_uart_1_avalon_jtag_slave_arb_share_counter_next_value assignment, which is an e_assign
  jtag_uart_1_avalon_jtag_slave_arb_share_counter_next_value <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(jtag_uart_1_avalon_jtag_slave_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(jtag_uart_1_avalon_jtag_slave_arb_share_set_values))) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(jtag_uart_1_avalon_jtag_slave_arb_share_counter) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(jtag_uart_1_avalon_jtag_slave_arb_share_counter))) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))));
  --jtag_uart_1_avalon_jtag_slave_allgrants all slave grants, which is an e_mux
  jtag_uart_1_avalon_jtag_slave_allgrants <= jtag_uart_1_avalon_jtag_slave_grant_vector;
  --jtag_uart_1_avalon_jtag_slave_end_xfer assignment, which is an e_assign
  jtag_uart_1_avalon_jtag_slave_end_xfer <= NOT ((jtag_uart_1_avalon_jtag_slave_waits_for_read OR jtag_uart_1_avalon_jtag_slave_waits_for_write));
  --end_xfer_arb_share_counter_term_jtag_uart_1_avalon_jtag_slave arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_jtag_uart_1_avalon_jtag_slave <= jtag_uart_1_avalon_jtag_slave_end_xfer AND (((NOT jtag_uart_1_avalon_jtag_slave_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --jtag_uart_1_avalon_jtag_slave_arb_share_counter arbitration counter enable, which is an e_assign
  jtag_uart_1_avalon_jtag_slave_arb_counter_enable <= ((end_xfer_arb_share_counter_term_jtag_uart_1_avalon_jtag_slave AND jtag_uart_1_avalon_jtag_slave_allgrants)) OR ((end_xfer_arb_share_counter_term_jtag_uart_1_avalon_jtag_slave AND NOT jtag_uart_1_avalon_jtag_slave_non_bursting_master_requests));
  --jtag_uart_1_avalon_jtag_slave_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      jtag_uart_1_avalon_jtag_slave_arb_share_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(jtag_uart_1_avalon_jtag_slave_arb_counter_enable) = '1' then 
        jtag_uart_1_avalon_jtag_slave_arb_share_counter <= jtag_uart_1_avalon_jtag_slave_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --jtag_uart_1_avalon_jtag_slave_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      jtag_uart_1_avalon_jtag_slave_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((jtag_uart_1_avalon_jtag_slave_master_qreq_vector AND end_xfer_arb_share_counter_term_jtag_uart_1_avalon_jtag_slave)) OR ((end_xfer_arb_share_counter_term_jtag_uart_1_avalon_jtag_slave AND NOT jtag_uart_1_avalon_jtag_slave_non_bursting_master_requests)))) = '1' then 
        jtag_uart_1_avalon_jtag_slave_slavearbiterlockenable <= jtag_uart_1_avalon_jtag_slave_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --ap_cpu/data_master jtag_uart_1/avalon_jtag_slave arbiterlock, which is an e_assign
  ap_cpu_data_master_arbiterlock <= jtag_uart_1_avalon_jtag_slave_slavearbiterlockenable AND ap_cpu_data_master_continuerequest;
  --jtag_uart_1_avalon_jtag_slave_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  jtag_uart_1_avalon_jtag_slave_slavearbiterlockenable2 <= jtag_uart_1_avalon_jtag_slave_arb_share_counter_next_value;
  --ap_cpu/data_master jtag_uart_1/avalon_jtag_slave arbiterlock2, which is an e_assign
  ap_cpu_data_master_arbiterlock2 <= jtag_uart_1_avalon_jtag_slave_slavearbiterlockenable2 AND ap_cpu_data_master_continuerequest;
  --jtag_uart_1_avalon_jtag_slave_any_continuerequest at least one master continues requesting, which is an e_assign
  jtag_uart_1_avalon_jtag_slave_any_continuerequest <= std_logic'('1');
  --ap_cpu_data_master_continuerequest continued request, which is an e_assign
  ap_cpu_data_master_continuerequest <= std_logic'('1');
  internal_ap_cpu_data_master_qualified_request_jtag_uart_1_avalon_jtag_slave <= internal_ap_cpu_data_master_requests_jtag_uart_1_avalon_jtag_slave AND NOT ((((ap_cpu_data_master_read AND (NOT ap_cpu_data_master_waitrequest))) OR (((NOT ap_cpu_data_master_waitrequest) AND ap_cpu_data_master_write))));
  --jtag_uart_1_avalon_jtag_slave_writedata mux, which is an e_mux
  jtag_uart_1_avalon_jtag_slave_writedata <= ap_cpu_data_master_writedata;
  --master is always granted when requested
  internal_ap_cpu_data_master_granted_jtag_uart_1_avalon_jtag_slave <= internal_ap_cpu_data_master_qualified_request_jtag_uart_1_avalon_jtag_slave;
  --ap_cpu/data_master saved-grant jtag_uart_1/avalon_jtag_slave, which is an e_assign
  ap_cpu_data_master_saved_grant_jtag_uart_1_avalon_jtag_slave <= internal_ap_cpu_data_master_requests_jtag_uart_1_avalon_jtag_slave;
  --allow new arb cycle for jtag_uart_1/avalon_jtag_slave, which is an e_assign
  jtag_uart_1_avalon_jtag_slave_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  jtag_uart_1_avalon_jtag_slave_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  jtag_uart_1_avalon_jtag_slave_master_qreq_vector <= std_logic'('1');
  --jtag_uart_1_avalon_jtag_slave_reset_n assignment, which is an e_assign
  jtag_uart_1_avalon_jtag_slave_reset_n <= reset_n;
  jtag_uart_1_avalon_jtag_slave_chipselect <= internal_ap_cpu_data_master_granted_jtag_uart_1_avalon_jtag_slave;
  --jtag_uart_1_avalon_jtag_slave_firsttransfer first transaction, which is an e_assign
  jtag_uart_1_avalon_jtag_slave_firsttransfer <= A_WE_StdLogic((std_logic'(jtag_uart_1_avalon_jtag_slave_begins_xfer) = '1'), jtag_uart_1_avalon_jtag_slave_unreg_firsttransfer, jtag_uart_1_avalon_jtag_slave_reg_firsttransfer);
  --jtag_uart_1_avalon_jtag_slave_unreg_firsttransfer first transaction, which is an e_assign
  jtag_uart_1_avalon_jtag_slave_unreg_firsttransfer <= NOT ((jtag_uart_1_avalon_jtag_slave_slavearbiterlockenable AND jtag_uart_1_avalon_jtag_slave_any_continuerequest));
  --jtag_uart_1_avalon_jtag_slave_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      jtag_uart_1_avalon_jtag_slave_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(jtag_uart_1_avalon_jtag_slave_begins_xfer) = '1' then 
        jtag_uart_1_avalon_jtag_slave_reg_firsttransfer <= jtag_uart_1_avalon_jtag_slave_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --jtag_uart_1_avalon_jtag_slave_beginbursttransfer_internal begin burst transfer, which is an e_assign
  jtag_uart_1_avalon_jtag_slave_beginbursttransfer_internal <= jtag_uart_1_avalon_jtag_slave_begins_xfer;
  --~jtag_uart_1_avalon_jtag_slave_read_n assignment, which is an e_mux
  jtag_uart_1_avalon_jtag_slave_read_n <= NOT ((internal_ap_cpu_data_master_granted_jtag_uart_1_avalon_jtag_slave AND ap_cpu_data_master_read));
  --~jtag_uart_1_avalon_jtag_slave_write_n assignment, which is an e_mux
  jtag_uart_1_avalon_jtag_slave_write_n <= NOT ((internal_ap_cpu_data_master_granted_jtag_uart_1_avalon_jtag_slave AND ap_cpu_data_master_write));
  shifted_address_to_jtag_uart_1_avalon_jtag_slave_from_ap_cpu_data_master <= ap_cpu_data_master_address_to_slave;
  --jtag_uart_1_avalon_jtag_slave_address mux, which is an e_mux
  jtag_uart_1_avalon_jtag_slave_address <= Vector_To_Std_Logic(A_SRL(shifted_address_to_jtag_uart_1_avalon_jtag_slave_from_ap_cpu_data_master,std_logic_vector'("00000000000000000000000000000010")));
  --d1_jtag_uart_1_avalon_jtag_slave_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_jtag_uart_1_avalon_jtag_slave_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_jtag_uart_1_avalon_jtag_slave_end_xfer <= jtag_uart_1_avalon_jtag_slave_end_xfer;
    end if;

  end process;

  --jtag_uart_1_avalon_jtag_slave_waits_for_read in a cycle, which is an e_mux
  jtag_uart_1_avalon_jtag_slave_waits_for_read <= jtag_uart_1_avalon_jtag_slave_in_a_read_cycle AND internal_jtag_uart_1_avalon_jtag_slave_waitrequest_from_sa;
  --jtag_uart_1_avalon_jtag_slave_in_a_read_cycle assignment, which is an e_assign
  jtag_uart_1_avalon_jtag_slave_in_a_read_cycle <= internal_ap_cpu_data_master_granted_jtag_uart_1_avalon_jtag_slave AND ap_cpu_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= jtag_uart_1_avalon_jtag_slave_in_a_read_cycle;
  --jtag_uart_1_avalon_jtag_slave_waits_for_write in a cycle, which is an e_mux
  jtag_uart_1_avalon_jtag_slave_waits_for_write <= jtag_uart_1_avalon_jtag_slave_in_a_write_cycle AND internal_jtag_uart_1_avalon_jtag_slave_waitrequest_from_sa;
  --jtag_uart_1_avalon_jtag_slave_in_a_write_cycle assignment, which is an e_assign
  jtag_uart_1_avalon_jtag_slave_in_a_write_cycle <= internal_ap_cpu_data_master_granted_jtag_uart_1_avalon_jtag_slave AND ap_cpu_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= jtag_uart_1_avalon_jtag_slave_in_a_write_cycle;
  wait_for_jtag_uart_1_avalon_jtag_slave_counter <= std_logic'('0');
  --assign jtag_uart_1_avalon_jtag_slave_irq_from_sa = jtag_uart_1_avalon_jtag_slave_irq so that symbol knows where to group signals which may go to master only, which is an e_assign
  jtag_uart_1_avalon_jtag_slave_irq_from_sa <= jtag_uart_1_avalon_jtag_slave_irq;
  --vhdl renameroo for output signals
  ap_cpu_data_master_granted_jtag_uart_1_avalon_jtag_slave <= internal_ap_cpu_data_master_granted_jtag_uart_1_avalon_jtag_slave;
  --vhdl renameroo for output signals
  ap_cpu_data_master_qualified_request_jtag_uart_1_avalon_jtag_slave <= internal_ap_cpu_data_master_qualified_request_jtag_uart_1_avalon_jtag_slave;
  --vhdl renameroo for output signals
  ap_cpu_data_master_requests_jtag_uart_1_avalon_jtag_slave <= internal_ap_cpu_data_master_requests_jtag_uart_1_avalon_jtag_slave;
  --vhdl renameroo for output signals
  jtag_uart_1_avalon_jtag_slave_waitrequest_from_sa <= internal_jtag_uart_1_avalon_jtag_slave_waitrequest_from_sa;
--synthesis translate_off
    --jtag_uart_1/avalon_jtag_slave enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity niosII_openMac_clock_0_in_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal niosII_openMac_clock_0_in_endofpacket : IN STD_LOGIC;
                 signal niosII_openMac_clock_0_in_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal niosII_openMac_clock_0_in_waitrequest : IN STD_LOGIC;
                 signal pcp_cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (25 DOWNTO 0);
                 signal pcp_cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal pcp_cpu_data_master_read : IN STD_LOGIC;
                 signal pcp_cpu_data_master_waitrequest : IN STD_LOGIC;
                 signal pcp_cpu_data_master_write : IN STD_LOGIC;
                 signal pcp_cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal d1_niosII_openMac_clock_0_in_end_xfer : OUT STD_LOGIC;
                 signal niosII_openMac_clock_0_in_address : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal niosII_openMac_clock_0_in_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal niosII_openMac_clock_0_in_endofpacket_from_sa : OUT STD_LOGIC;
                 signal niosII_openMac_clock_0_in_nativeaddress : OUT STD_LOGIC;
                 signal niosII_openMac_clock_0_in_read : OUT STD_LOGIC;
                 signal niosII_openMac_clock_0_in_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal niosII_openMac_clock_0_in_reset_n : OUT STD_LOGIC;
                 signal niosII_openMac_clock_0_in_waitrequest_from_sa : OUT STD_LOGIC;
                 signal niosII_openMac_clock_0_in_write : OUT STD_LOGIC;
                 signal niosII_openMac_clock_0_in_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal pcp_cpu_data_master_granted_niosII_openMac_clock_0_in : OUT STD_LOGIC;
                 signal pcp_cpu_data_master_qualified_request_niosII_openMac_clock_0_in : OUT STD_LOGIC;
                 signal pcp_cpu_data_master_read_data_valid_niosII_openMac_clock_0_in : OUT STD_LOGIC;
                 signal pcp_cpu_data_master_requests_niosII_openMac_clock_0_in : OUT STD_LOGIC
              );
end entity niosII_openMac_clock_0_in_arbitrator;


architecture europa of niosII_openMac_clock_0_in_arbitrator is
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_niosII_openMac_clock_0_in :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_niosII_openMac_clock_0_in_waitrequest_from_sa :  STD_LOGIC;
                signal internal_pcp_cpu_data_master_granted_niosII_openMac_clock_0_in :  STD_LOGIC;
                signal internal_pcp_cpu_data_master_qualified_request_niosII_openMac_clock_0_in :  STD_LOGIC;
                signal internal_pcp_cpu_data_master_requests_niosII_openMac_clock_0_in :  STD_LOGIC;
                signal niosII_openMac_clock_0_in_allgrants :  STD_LOGIC;
                signal niosII_openMac_clock_0_in_allow_new_arb_cycle :  STD_LOGIC;
                signal niosII_openMac_clock_0_in_any_bursting_master_saved_grant :  STD_LOGIC;
                signal niosII_openMac_clock_0_in_any_continuerequest :  STD_LOGIC;
                signal niosII_openMac_clock_0_in_arb_counter_enable :  STD_LOGIC;
                signal niosII_openMac_clock_0_in_arb_share_counter :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal niosII_openMac_clock_0_in_arb_share_counter_next_value :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal niosII_openMac_clock_0_in_arb_share_set_values :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal niosII_openMac_clock_0_in_beginbursttransfer_internal :  STD_LOGIC;
                signal niosII_openMac_clock_0_in_begins_xfer :  STD_LOGIC;
                signal niosII_openMac_clock_0_in_end_xfer :  STD_LOGIC;
                signal niosII_openMac_clock_0_in_firsttransfer :  STD_LOGIC;
                signal niosII_openMac_clock_0_in_grant_vector :  STD_LOGIC;
                signal niosII_openMac_clock_0_in_in_a_read_cycle :  STD_LOGIC;
                signal niosII_openMac_clock_0_in_in_a_write_cycle :  STD_LOGIC;
                signal niosII_openMac_clock_0_in_master_qreq_vector :  STD_LOGIC;
                signal niosII_openMac_clock_0_in_non_bursting_master_requests :  STD_LOGIC;
                signal niosII_openMac_clock_0_in_reg_firsttransfer :  STD_LOGIC;
                signal niosII_openMac_clock_0_in_slavearbiterlockenable :  STD_LOGIC;
                signal niosII_openMac_clock_0_in_slavearbiterlockenable2 :  STD_LOGIC;
                signal niosII_openMac_clock_0_in_unreg_firsttransfer :  STD_LOGIC;
                signal niosII_openMac_clock_0_in_waits_for_read :  STD_LOGIC;
                signal niosII_openMac_clock_0_in_waits_for_write :  STD_LOGIC;
                signal pcp_cpu_data_master_arbiterlock :  STD_LOGIC;
                signal pcp_cpu_data_master_arbiterlock2 :  STD_LOGIC;
                signal pcp_cpu_data_master_continuerequest :  STD_LOGIC;
                signal pcp_cpu_data_master_saved_grant_niosII_openMac_clock_0_in :  STD_LOGIC;
                signal shifted_address_to_niosII_openMac_clock_0_in_from_pcp_cpu_data_master :  STD_LOGIC_VECTOR (25 DOWNTO 0);
                signal wait_for_niosII_openMac_clock_0_in_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT niosII_openMac_clock_0_in_end_xfer;
    end if;

  end process;

  niosII_openMac_clock_0_in_begins_xfer <= NOT d1_reasons_to_wait AND (internal_pcp_cpu_data_master_qualified_request_niosII_openMac_clock_0_in);
  --assign niosII_openMac_clock_0_in_readdata_from_sa = niosII_openMac_clock_0_in_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  niosII_openMac_clock_0_in_readdata_from_sa <= niosII_openMac_clock_0_in_readdata;
  internal_pcp_cpu_data_master_requests_niosII_openMac_clock_0_in <= to_std_logic(((Std_Logic_Vector'(pcp_cpu_data_master_address_to_slave(25 DOWNTO 3) & std_logic_vector'("000")) = std_logic_vector'("00000000000000100100011000")))) AND ((pcp_cpu_data_master_read OR pcp_cpu_data_master_write));
  --assign niosII_openMac_clock_0_in_waitrequest_from_sa = niosII_openMac_clock_0_in_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_niosII_openMac_clock_0_in_waitrequest_from_sa <= niosII_openMac_clock_0_in_waitrequest;
  --niosII_openMac_clock_0_in_arb_share_counter set values, which is an e_mux
  niosII_openMac_clock_0_in_arb_share_set_values <= std_logic_vector'("01");
  --niosII_openMac_clock_0_in_non_bursting_master_requests mux, which is an e_mux
  niosII_openMac_clock_0_in_non_bursting_master_requests <= internal_pcp_cpu_data_master_requests_niosII_openMac_clock_0_in;
  --niosII_openMac_clock_0_in_any_bursting_master_saved_grant mux, which is an e_mux
  niosII_openMac_clock_0_in_any_bursting_master_saved_grant <= std_logic'('0');
  --niosII_openMac_clock_0_in_arb_share_counter_next_value assignment, which is an e_assign
  niosII_openMac_clock_0_in_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(niosII_openMac_clock_0_in_firsttransfer) = '1'), (((std_logic_vector'("0000000000000000000000000000000") & (niosII_openMac_clock_0_in_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(niosII_openMac_clock_0_in_arb_share_counter)) = '1'), (((std_logic_vector'("0000000000000000000000000000000") & (niosII_openMac_clock_0_in_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 2);
  --niosII_openMac_clock_0_in_allgrants all slave grants, which is an e_mux
  niosII_openMac_clock_0_in_allgrants <= niosII_openMac_clock_0_in_grant_vector;
  --niosII_openMac_clock_0_in_end_xfer assignment, which is an e_assign
  niosII_openMac_clock_0_in_end_xfer <= NOT ((niosII_openMac_clock_0_in_waits_for_read OR niosII_openMac_clock_0_in_waits_for_write));
  --end_xfer_arb_share_counter_term_niosII_openMac_clock_0_in arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_niosII_openMac_clock_0_in <= niosII_openMac_clock_0_in_end_xfer AND (((NOT niosII_openMac_clock_0_in_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --niosII_openMac_clock_0_in_arb_share_counter arbitration counter enable, which is an e_assign
  niosII_openMac_clock_0_in_arb_counter_enable <= ((end_xfer_arb_share_counter_term_niosII_openMac_clock_0_in AND niosII_openMac_clock_0_in_allgrants)) OR ((end_xfer_arb_share_counter_term_niosII_openMac_clock_0_in AND NOT niosII_openMac_clock_0_in_non_bursting_master_requests));
  --niosII_openMac_clock_0_in_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_openMac_clock_0_in_arb_share_counter <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      if std_logic'(niosII_openMac_clock_0_in_arb_counter_enable) = '1' then 
        niosII_openMac_clock_0_in_arb_share_counter <= niosII_openMac_clock_0_in_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --niosII_openMac_clock_0_in_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_openMac_clock_0_in_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((niosII_openMac_clock_0_in_master_qreq_vector AND end_xfer_arb_share_counter_term_niosII_openMac_clock_0_in)) OR ((end_xfer_arb_share_counter_term_niosII_openMac_clock_0_in AND NOT niosII_openMac_clock_0_in_non_bursting_master_requests)))) = '1' then 
        niosII_openMac_clock_0_in_slavearbiterlockenable <= or_reduce(niosII_openMac_clock_0_in_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --pcp_cpu/data_master niosII_openMac_clock_0/in arbiterlock, which is an e_assign
  pcp_cpu_data_master_arbiterlock <= niosII_openMac_clock_0_in_slavearbiterlockenable AND pcp_cpu_data_master_continuerequest;
  --niosII_openMac_clock_0_in_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  niosII_openMac_clock_0_in_slavearbiterlockenable2 <= or_reduce(niosII_openMac_clock_0_in_arb_share_counter_next_value);
  --pcp_cpu/data_master niosII_openMac_clock_0/in arbiterlock2, which is an e_assign
  pcp_cpu_data_master_arbiterlock2 <= niosII_openMac_clock_0_in_slavearbiterlockenable2 AND pcp_cpu_data_master_continuerequest;
  --niosII_openMac_clock_0_in_any_continuerequest at least one master continues requesting, which is an e_assign
  niosII_openMac_clock_0_in_any_continuerequest <= std_logic'('1');
  --pcp_cpu_data_master_continuerequest continued request, which is an e_assign
  pcp_cpu_data_master_continuerequest <= std_logic'('1');
  internal_pcp_cpu_data_master_qualified_request_niosII_openMac_clock_0_in <= internal_pcp_cpu_data_master_requests_niosII_openMac_clock_0_in AND NOT ((((pcp_cpu_data_master_read AND (NOT pcp_cpu_data_master_waitrequest))) OR (((NOT pcp_cpu_data_master_waitrequest) AND pcp_cpu_data_master_write))));
  --niosII_openMac_clock_0_in_writedata mux, which is an e_mux
  niosII_openMac_clock_0_in_writedata <= pcp_cpu_data_master_writedata;
  --assign niosII_openMac_clock_0_in_endofpacket_from_sa = niosII_openMac_clock_0_in_endofpacket so that symbol knows where to group signals which may go to master only, which is an e_assign
  niosII_openMac_clock_0_in_endofpacket_from_sa <= niosII_openMac_clock_0_in_endofpacket;
  --master is always granted when requested
  internal_pcp_cpu_data_master_granted_niosII_openMac_clock_0_in <= internal_pcp_cpu_data_master_qualified_request_niosII_openMac_clock_0_in;
  --pcp_cpu/data_master saved-grant niosII_openMac_clock_0/in, which is an e_assign
  pcp_cpu_data_master_saved_grant_niosII_openMac_clock_0_in <= internal_pcp_cpu_data_master_requests_niosII_openMac_clock_0_in;
  --allow new arb cycle for niosII_openMac_clock_0/in, which is an e_assign
  niosII_openMac_clock_0_in_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  niosII_openMac_clock_0_in_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  niosII_openMac_clock_0_in_master_qreq_vector <= std_logic'('1');
  --niosII_openMac_clock_0_in_reset_n assignment, which is an e_assign
  niosII_openMac_clock_0_in_reset_n <= reset_n;
  --niosII_openMac_clock_0_in_firsttransfer first transaction, which is an e_assign
  niosII_openMac_clock_0_in_firsttransfer <= A_WE_StdLogic((std_logic'(niosII_openMac_clock_0_in_begins_xfer) = '1'), niosII_openMac_clock_0_in_unreg_firsttransfer, niosII_openMac_clock_0_in_reg_firsttransfer);
  --niosII_openMac_clock_0_in_unreg_firsttransfer first transaction, which is an e_assign
  niosII_openMac_clock_0_in_unreg_firsttransfer <= NOT ((niosII_openMac_clock_0_in_slavearbiterlockenable AND niosII_openMac_clock_0_in_any_continuerequest));
  --niosII_openMac_clock_0_in_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_openMac_clock_0_in_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(niosII_openMac_clock_0_in_begins_xfer) = '1' then 
        niosII_openMac_clock_0_in_reg_firsttransfer <= niosII_openMac_clock_0_in_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --niosII_openMac_clock_0_in_beginbursttransfer_internal begin burst transfer, which is an e_assign
  niosII_openMac_clock_0_in_beginbursttransfer_internal <= niosII_openMac_clock_0_in_begins_xfer;
  --niosII_openMac_clock_0_in_read assignment, which is an e_mux
  niosII_openMac_clock_0_in_read <= internal_pcp_cpu_data_master_granted_niosII_openMac_clock_0_in AND pcp_cpu_data_master_read;
  --niosII_openMac_clock_0_in_write assignment, which is an e_mux
  niosII_openMac_clock_0_in_write <= internal_pcp_cpu_data_master_granted_niosII_openMac_clock_0_in AND pcp_cpu_data_master_write;
  shifted_address_to_niosII_openMac_clock_0_in_from_pcp_cpu_data_master <= pcp_cpu_data_master_address_to_slave;
  --niosII_openMac_clock_0_in_address mux, which is an e_mux
  niosII_openMac_clock_0_in_address <= A_EXT (A_SRL(shifted_address_to_niosII_openMac_clock_0_in_from_pcp_cpu_data_master,std_logic_vector'("00000000000000000000000000000010")), 3);
  --slaveid niosII_openMac_clock_0_in_nativeaddress nativeaddress mux, which is an e_mux
  niosII_openMac_clock_0_in_nativeaddress <= Vector_To_Std_Logic(A_SRL(pcp_cpu_data_master_address_to_slave,std_logic_vector'("00000000000000000000000000000010")));
  --d1_niosII_openMac_clock_0_in_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_niosII_openMac_clock_0_in_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_niosII_openMac_clock_0_in_end_xfer <= niosII_openMac_clock_0_in_end_xfer;
    end if;

  end process;

  --niosII_openMac_clock_0_in_waits_for_read in a cycle, which is an e_mux
  niosII_openMac_clock_0_in_waits_for_read <= niosII_openMac_clock_0_in_in_a_read_cycle AND internal_niosII_openMac_clock_0_in_waitrequest_from_sa;
  --niosII_openMac_clock_0_in_in_a_read_cycle assignment, which is an e_assign
  niosII_openMac_clock_0_in_in_a_read_cycle <= internal_pcp_cpu_data_master_granted_niosII_openMac_clock_0_in AND pcp_cpu_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= niosII_openMac_clock_0_in_in_a_read_cycle;
  --niosII_openMac_clock_0_in_waits_for_write in a cycle, which is an e_mux
  niosII_openMac_clock_0_in_waits_for_write <= niosII_openMac_clock_0_in_in_a_write_cycle AND internal_niosII_openMac_clock_0_in_waitrequest_from_sa;
  --niosII_openMac_clock_0_in_in_a_write_cycle assignment, which is an e_assign
  niosII_openMac_clock_0_in_in_a_write_cycle <= internal_pcp_cpu_data_master_granted_niosII_openMac_clock_0_in AND pcp_cpu_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= niosII_openMac_clock_0_in_in_a_write_cycle;
  wait_for_niosII_openMac_clock_0_in_counter <= std_logic'('0');
  --niosII_openMac_clock_0_in_byteenable byte enable port mux, which is an e_mux
  niosII_openMac_clock_0_in_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_pcp_cpu_data_master_granted_niosII_openMac_clock_0_in)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (pcp_cpu_data_master_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))), 4);
  --vhdl renameroo for output signals
  niosII_openMac_clock_0_in_waitrequest_from_sa <= internal_niosII_openMac_clock_0_in_waitrequest_from_sa;
  --vhdl renameroo for output signals
  pcp_cpu_data_master_granted_niosII_openMac_clock_0_in <= internal_pcp_cpu_data_master_granted_niosII_openMac_clock_0_in;
  --vhdl renameroo for output signals
  pcp_cpu_data_master_qualified_request_niosII_openMac_clock_0_in <= internal_pcp_cpu_data_master_qualified_request_niosII_openMac_clock_0_in;
  --vhdl renameroo for output signals
  pcp_cpu_data_master_requests_niosII_openMac_clock_0_in <= internal_pcp_cpu_data_master_requests_niosII_openMac_clock_0_in;
--synthesis translate_off
    --niosII_openMac_clock_0/in enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity niosII_openMac_clock_0_out_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal d1_jtag_uart_0_avalon_jtag_slave_end_xfer : IN STD_LOGIC;
                 signal jtag_uart_0_avalon_jtag_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal jtag_uart_0_avalon_jtag_slave_waitrequest_from_sa : IN STD_LOGIC;
                 signal niosII_openMac_clock_0_out_address : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal niosII_openMac_clock_0_out_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal niosII_openMac_clock_0_out_granted_jtag_uart_0_avalon_jtag_slave : IN STD_LOGIC;
                 signal niosII_openMac_clock_0_out_qualified_request_jtag_uart_0_avalon_jtag_slave : IN STD_LOGIC;
                 signal niosII_openMac_clock_0_out_read : IN STD_LOGIC;
                 signal niosII_openMac_clock_0_out_read_data_valid_jtag_uart_0_avalon_jtag_slave : IN STD_LOGIC;
                 signal niosII_openMac_clock_0_out_requests_jtag_uart_0_avalon_jtag_slave : IN STD_LOGIC;
                 signal niosII_openMac_clock_0_out_write : IN STD_LOGIC;
                 signal niosII_openMac_clock_0_out_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal niosII_openMac_clock_0_out_address_to_slave : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal niosII_openMac_clock_0_out_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal niosII_openMac_clock_0_out_reset_n : OUT STD_LOGIC;
                 signal niosII_openMac_clock_0_out_waitrequest : OUT STD_LOGIC
              );
end entity niosII_openMac_clock_0_out_arbitrator;


architecture europa of niosII_openMac_clock_0_out_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal internal_niosII_openMac_clock_0_out_address_to_slave :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal internal_niosII_openMac_clock_0_out_waitrequest :  STD_LOGIC;
                signal niosII_openMac_clock_0_out_address_last_time :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal niosII_openMac_clock_0_out_byteenable_last_time :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_openMac_clock_0_out_read_last_time :  STD_LOGIC;
                signal niosII_openMac_clock_0_out_run :  STD_LOGIC;
                signal niosII_openMac_clock_0_out_write_last_time :  STD_LOGIC;
                signal niosII_openMac_clock_0_out_writedata_last_time :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal r_0 :  STD_LOGIC;

begin

  --r_0 master_run cascaded wait assignment, which is an e_assign
  r_0 <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000001") AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT niosII_openMac_clock_0_out_qualified_request_jtag_uart_0_avalon_jtag_slave OR NOT ((niosII_openMac_clock_0_out_read OR niosII_openMac_clock_0_out_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT jtag_uart_0_avalon_jtag_slave_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((niosII_openMac_clock_0_out_read OR niosII_openMac_clock_0_out_write)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT niosII_openMac_clock_0_out_qualified_request_jtag_uart_0_avalon_jtag_slave OR NOT ((niosII_openMac_clock_0_out_read OR niosII_openMac_clock_0_out_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT jtag_uart_0_avalon_jtag_slave_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((niosII_openMac_clock_0_out_read OR niosII_openMac_clock_0_out_write)))))))))));
  --cascaded wait assignment, which is an e_assign
  niosII_openMac_clock_0_out_run <= r_0;
  --optimize select-logic by passing only those address bits which matter.
  internal_niosII_openMac_clock_0_out_address_to_slave <= niosII_openMac_clock_0_out_address;
  --niosII_openMac_clock_0/out readdata mux, which is an e_mux
  niosII_openMac_clock_0_out_readdata <= jtag_uart_0_avalon_jtag_slave_readdata_from_sa;
  --actual waitrequest port, which is an e_assign
  internal_niosII_openMac_clock_0_out_waitrequest <= NOT niosII_openMac_clock_0_out_run;
  --niosII_openMac_clock_0_out_reset_n assignment, which is an e_assign
  niosII_openMac_clock_0_out_reset_n <= reset_n;
  --vhdl renameroo for output signals
  niosII_openMac_clock_0_out_address_to_slave <= internal_niosII_openMac_clock_0_out_address_to_slave;
  --vhdl renameroo for output signals
  niosII_openMac_clock_0_out_waitrequest <= internal_niosII_openMac_clock_0_out_waitrequest;
--synthesis translate_off
    --niosII_openMac_clock_0_out_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_openMac_clock_0_out_address_last_time <= std_logic_vector'("000");
      elsif clk'event and clk = '1' then
        niosII_openMac_clock_0_out_address_last_time <= niosII_openMac_clock_0_out_address;
      end if;

    end process;

    --niosII_openMac_clock_0/out waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_niosII_openMac_clock_0_out_waitrequest AND ((niosII_openMac_clock_0_out_read OR niosII_openMac_clock_0_out_write));
      end if;

    end process;

    --niosII_openMac_clock_0_out_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line16 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((niosII_openMac_clock_0_out_address /= niosII_openMac_clock_0_out_address_last_time))))) = '1' then 
          write(write_line16, now);
          write(write_line16, string'(": "));
          write(write_line16, string'("niosII_openMac_clock_0_out_address did not heed wait!!!"));
          write(output, write_line16.all);
          deallocate (write_line16);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_openMac_clock_0_out_byteenable check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_openMac_clock_0_out_byteenable_last_time <= std_logic_vector'("0000");
      elsif clk'event and clk = '1' then
        niosII_openMac_clock_0_out_byteenable_last_time <= niosII_openMac_clock_0_out_byteenable;
      end if;

    end process;

    --niosII_openMac_clock_0_out_byteenable matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line17 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((niosII_openMac_clock_0_out_byteenable /= niosII_openMac_clock_0_out_byteenable_last_time))))) = '1' then 
          write(write_line17, now);
          write(write_line17, string'(": "));
          write(write_line17, string'("niosII_openMac_clock_0_out_byteenable did not heed wait!!!"));
          write(output, write_line17.all);
          deallocate (write_line17);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_openMac_clock_0_out_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_openMac_clock_0_out_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        niosII_openMac_clock_0_out_read_last_time <= niosII_openMac_clock_0_out_read;
      end if;

    end process;

    --niosII_openMac_clock_0_out_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line18 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(niosII_openMac_clock_0_out_read) /= std_logic'(niosII_openMac_clock_0_out_read_last_time)))))) = '1' then 
          write(write_line18, now);
          write(write_line18, string'(": "));
          write(write_line18, string'("niosII_openMac_clock_0_out_read did not heed wait!!!"));
          write(output, write_line18.all);
          deallocate (write_line18);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_openMac_clock_0_out_write check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_openMac_clock_0_out_write_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        niosII_openMac_clock_0_out_write_last_time <= niosII_openMac_clock_0_out_write;
      end if;

    end process;

    --niosII_openMac_clock_0_out_write matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line19 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(niosII_openMac_clock_0_out_write) /= std_logic'(niosII_openMac_clock_0_out_write_last_time)))))) = '1' then 
          write(write_line19, now);
          write(write_line19, string'(": "));
          write(write_line19, string'("niosII_openMac_clock_0_out_write did not heed wait!!!"));
          write(output, write_line19.all);
          deallocate (write_line19);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_openMac_clock_0_out_writedata check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_openMac_clock_0_out_writedata_last_time <= std_logic_vector'("00000000000000000000000000000000");
      elsif clk'event and clk = '1' then
        niosII_openMac_clock_0_out_writedata_last_time <= niosII_openMac_clock_0_out_writedata;
      end if;

    end process;

    --niosII_openMac_clock_0_out_writedata matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line20 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((active_and_waiting_last_time AND to_std_logic(((niosII_openMac_clock_0_out_writedata /= niosII_openMac_clock_0_out_writedata_last_time)))) AND niosII_openMac_clock_0_out_write)) = '1' then 
          write(write_line20, now);
          write(write_line20, string'(": "));
          write(write_line20, string'("niosII_openMac_clock_0_out_writedata did not heed wait!!!"));
          write(output, write_line20.all);
          deallocate (write_line20);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity niosII_openMac_clock_1_in_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal niosII_openMac_clock_1_in_endofpacket : IN STD_LOGIC;
                 signal niosII_openMac_clock_1_in_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal niosII_openMac_clock_1_in_waitrequest : IN STD_LOGIC;
                 signal pcp_cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (25 DOWNTO 0);
                 signal pcp_cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal pcp_cpu_data_master_read : IN STD_LOGIC;
                 signal pcp_cpu_data_master_waitrequest : IN STD_LOGIC;
                 signal pcp_cpu_data_master_write : IN STD_LOGIC;
                 signal pcp_cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal d1_niosII_openMac_clock_1_in_end_xfer : OUT STD_LOGIC;
                 signal niosII_openMac_clock_1_in_address : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal niosII_openMac_clock_1_in_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal niosII_openMac_clock_1_in_endofpacket_from_sa : OUT STD_LOGIC;
                 signal niosII_openMac_clock_1_in_nativeaddress : OUT STD_LOGIC;
                 signal niosII_openMac_clock_1_in_read : OUT STD_LOGIC;
                 signal niosII_openMac_clock_1_in_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal niosII_openMac_clock_1_in_reset_n : OUT STD_LOGIC;
                 signal niosII_openMac_clock_1_in_waitrequest_from_sa : OUT STD_LOGIC;
                 signal niosII_openMac_clock_1_in_write : OUT STD_LOGIC;
                 signal niosII_openMac_clock_1_in_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal pcp_cpu_data_master_granted_niosII_openMac_clock_1_in : OUT STD_LOGIC;
                 signal pcp_cpu_data_master_qualified_request_niosII_openMac_clock_1_in : OUT STD_LOGIC;
                 signal pcp_cpu_data_master_read_data_valid_niosII_openMac_clock_1_in : OUT STD_LOGIC;
                 signal pcp_cpu_data_master_requests_niosII_openMac_clock_1_in : OUT STD_LOGIC
              );
end entity niosII_openMac_clock_1_in_arbitrator;


architecture europa of niosII_openMac_clock_1_in_arbitrator is
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_niosII_openMac_clock_1_in :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_niosII_openMac_clock_1_in_waitrequest_from_sa :  STD_LOGIC;
                signal internal_pcp_cpu_data_master_granted_niosII_openMac_clock_1_in :  STD_LOGIC;
                signal internal_pcp_cpu_data_master_qualified_request_niosII_openMac_clock_1_in :  STD_LOGIC;
                signal internal_pcp_cpu_data_master_requests_niosII_openMac_clock_1_in :  STD_LOGIC;
                signal niosII_openMac_clock_1_in_allgrants :  STD_LOGIC;
                signal niosII_openMac_clock_1_in_allow_new_arb_cycle :  STD_LOGIC;
                signal niosII_openMac_clock_1_in_any_bursting_master_saved_grant :  STD_LOGIC;
                signal niosII_openMac_clock_1_in_any_continuerequest :  STD_LOGIC;
                signal niosII_openMac_clock_1_in_arb_counter_enable :  STD_LOGIC;
                signal niosII_openMac_clock_1_in_arb_share_counter :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal niosII_openMac_clock_1_in_arb_share_counter_next_value :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal niosII_openMac_clock_1_in_arb_share_set_values :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal niosII_openMac_clock_1_in_beginbursttransfer_internal :  STD_LOGIC;
                signal niosII_openMac_clock_1_in_begins_xfer :  STD_LOGIC;
                signal niosII_openMac_clock_1_in_end_xfer :  STD_LOGIC;
                signal niosII_openMac_clock_1_in_firsttransfer :  STD_LOGIC;
                signal niosII_openMac_clock_1_in_grant_vector :  STD_LOGIC;
                signal niosII_openMac_clock_1_in_in_a_read_cycle :  STD_LOGIC;
                signal niosII_openMac_clock_1_in_in_a_write_cycle :  STD_LOGIC;
                signal niosII_openMac_clock_1_in_master_qreq_vector :  STD_LOGIC;
                signal niosII_openMac_clock_1_in_non_bursting_master_requests :  STD_LOGIC;
                signal niosII_openMac_clock_1_in_reg_firsttransfer :  STD_LOGIC;
                signal niosII_openMac_clock_1_in_slavearbiterlockenable :  STD_LOGIC;
                signal niosII_openMac_clock_1_in_slavearbiterlockenable2 :  STD_LOGIC;
                signal niosII_openMac_clock_1_in_unreg_firsttransfer :  STD_LOGIC;
                signal niosII_openMac_clock_1_in_waits_for_read :  STD_LOGIC;
                signal niosII_openMac_clock_1_in_waits_for_write :  STD_LOGIC;
                signal pcp_cpu_data_master_arbiterlock :  STD_LOGIC;
                signal pcp_cpu_data_master_arbiterlock2 :  STD_LOGIC;
                signal pcp_cpu_data_master_continuerequest :  STD_LOGIC;
                signal pcp_cpu_data_master_saved_grant_niosII_openMac_clock_1_in :  STD_LOGIC;
                signal wait_for_niosII_openMac_clock_1_in_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT niosII_openMac_clock_1_in_end_xfer;
    end if;

  end process;

  niosII_openMac_clock_1_in_begins_xfer <= NOT d1_reasons_to_wait AND (internal_pcp_cpu_data_master_qualified_request_niosII_openMac_clock_1_in);
  --assign niosII_openMac_clock_1_in_readdata_from_sa = niosII_openMac_clock_1_in_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  niosII_openMac_clock_1_in_readdata_from_sa <= niosII_openMac_clock_1_in_readdata;
  internal_pcp_cpu_data_master_requests_niosII_openMac_clock_1_in <= to_std_logic(((Std_Logic_Vector'(pcp_cpu_data_master_address_to_slave(25 DOWNTO 3) & std_logic_vector'("000")) = std_logic_vector'("00000000000000100100010000")))) AND ((pcp_cpu_data_master_read OR pcp_cpu_data_master_write));
  --assign niosII_openMac_clock_1_in_waitrequest_from_sa = niosII_openMac_clock_1_in_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_niosII_openMac_clock_1_in_waitrequest_from_sa <= niosII_openMac_clock_1_in_waitrequest;
  --niosII_openMac_clock_1_in_arb_share_counter set values, which is an e_mux
  niosII_openMac_clock_1_in_arb_share_set_values <= std_logic_vector'("01");
  --niosII_openMac_clock_1_in_non_bursting_master_requests mux, which is an e_mux
  niosII_openMac_clock_1_in_non_bursting_master_requests <= internal_pcp_cpu_data_master_requests_niosII_openMac_clock_1_in;
  --niosII_openMac_clock_1_in_any_bursting_master_saved_grant mux, which is an e_mux
  niosII_openMac_clock_1_in_any_bursting_master_saved_grant <= std_logic'('0');
  --niosII_openMac_clock_1_in_arb_share_counter_next_value assignment, which is an e_assign
  niosII_openMac_clock_1_in_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(niosII_openMac_clock_1_in_firsttransfer) = '1'), (((std_logic_vector'("0000000000000000000000000000000") & (niosII_openMac_clock_1_in_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(niosII_openMac_clock_1_in_arb_share_counter)) = '1'), (((std_logic_vector'("0000000000000000000000000000000") & (niosII_openMac_clock_1_in_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 2);
  --niosII_openMac_clock_1_in_allgrants all slave grants, which is an e_mux
  niosII_openMac_clock_1_in_allgrants <= niosII_openMac_clock_1_in_grant_vector;
  --niosII_openMac_clock_1_in_end_xfer assignment, which is an e_assign
  niosII_openMac_clock_1_in_end_xfer <= NOT ((niosII_openMac_clock_1_in_waits_for_read OR niosII_openMac_clock_1_in_waits_for_write));
  --end_xfer_arb_share_counter_term_niosII_openMac_clock_1_in arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_niosII_openMac_clock_1_in <= niosII_openMac_clock_1_in_end_xfer AND (((NOT niosII_openMac_clock_1_in_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --niosII_openMac_clock_1_in_arb_share_counter arbitration counter enable, which is an e_assign
  niosII_openMac_clock_1_in_arb_counter_enable <= ((end_xfer_arb_share_counter_term_niosII_openMac_clock_1_in AND niosII_openMac_clock_1_in_allgrants)) OR ((end_xfer_arb_share_counter_term_niosII_openMac_clock_1_in AND NOT niosII_openMac_clock_1_in_non_bursting_master_requests));
  --niosII_openMac_clock_1_in_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_openMac_clock_1_in_arb_share_counter <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      if std_logic'(niosII_openMac_clock_1_in_arb_counter_enable) = '1' then 
        niosII_openMac_clock_1_in_arb_share_counter <= niosII_openMac_clock_1_in_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --niosII_openMac_clock_1_in_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_openMac_clock_1_in_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((niosII_openMac_clock_1_in_master_qreq_vector AND end_xfer_arb_share_counter_term_niosII_openMac_clock_1_in)) OR ((end_xfer_arb_share_counter_term_niosII_openMac_clock_1_in AND NOT niosII_openMac_clock_1_in_non_bursting_master_requests)))) = '1' then 
        niosII_openMac_clock_1_in_slavearbiterlockenable <= or_reduce(niosII_openMac_clock_1_in_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --pcp_cpu/data_master niosII_openMac_clock_1/in arbiterlock, which is an e_assign
  pcp_cpu_data_master_arbiterlock <= niosII_openMac_clock_1_in_slavearbiterlockenable AND pcp_cpu_data_master_continuerequest;
  --niosII_openMac_clock_1_in_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  niosII_openMac_clock_1_in_slavearbiterlockenable2 <= or_reduce(niosII_openMac_clock_1_in_arb_share_counter_next_value);
  --pcp_cpu/data_master niosII_openMac_clock_1/in arbiterlock2, which is an e_assign
  pcp_cpu_data_master_arbiterlock2 <= niosII_openMac_clock_1_in_slavearbiterlockenable2 AND pcp_cpu_data_master_continuerequest;
  --niosII_openMac_clock_1_in_any_continuerequest at least one master continues requesting, which is an e_assign
  niosII_openMac_clock_1_in_any_continuerequest <= std_logic'('1');
  --pcp_cpu_data_master_continuerequest continued request, which is an e_assign
  pcp_cpu_data_master_continuerequest <= std_logic'('1');
  internal_pcp_cpu_data_master_qualified_request_niosII_openMac_clock_1_in <= internal_pcp_cpu_data_master_requests_niosII_openMac_clock_1_in AND NOT ((((pcp_cpu_data_master_read AND (NOT pcp_cpu_data_master_waitrequest))) OR (((NOT pcp_cpu_data_master_waitrequest) AND pcp_cpu_data_master_write))));
  --niosII_openMac_clock_1_in_writedata mux, which is an e_mux
  niosII_openMac_clock_1_in_writedata <= pcp_cpu_data_master_writedata;
  --assign niosII_openMac_clock_1_in_endofpacket_from_sa = niosII_openMac_clock_1_in_endofpacket so that symbol knows where to group signals which may go to master only, which is an e_assign
  niosII_openMac_clock_1_in_endofpacket_from_sa <= niosII_openMac_clock_1_in_endofpacket;
  --master is always granted when requested
  internal_pcp_cpu_data_master_granted_niosII_openMac_clock_1_in <= internal_pcp_cpu_data_master_qualified_request_niosII_openMac_clock_1_in;
  --pcp_cpu/data_master saved-grant niosII_openMac_clock_1/in, which is an e_assign
  pcp_cpu_data_master_saved_grant_niosII_openMac_clock_1_in <= internal_pcp_cpu_data_master_requests_niosII_openMac_clock_1_in;
  --allow new arb cycle for niosII_openMac_clock_1/in, which is an e_assign
  niosII_openMac_clock_1_in_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  niosII_openMac_clock_1_in_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  niosII_openMac_clock_1_in_master_qreq_vector <= std_logic'('1');
  --niosII_openMac_clock_1_in_reset_n assignment, which is an e_assign
  niosII_openMac_clock_1_in_reset_n <= reset_n;
  --niosII_openMac_clock_1_in_firsttransfer first transaction, which is an e_assign
  niosII_openMac_clock_1_in_firsttransfer <= A_WE_StdLogic((std_logic'(niosII_openMac_clock_1_in_begins_xfer) = '1'), niosII_openMac_clock_1_in_unreg_firsttransfer, niosII_openMac_clock_1_in_reg_firsttransfer);
  --niosII_openMac_clock_1_in_unreg_firsttransfer first transaction, which is an e_assign
  niosII_openMac_clock_1_in_unreg_firsttransfer <= NOT ((niosII_openMac_clock_1_in_slavearbiterlockenable AND niosII_openMac_clock_1_in_any_continuerequest));
  --niosII_openMac_clock_1_in_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_openMac_clock_1_in_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(niosII_openMac_clock_1_in_begins_xfer) = '1' then 
        niosII_openMac_clock_1_in_reg_firsttransfer <= niosII_openMac_clock_1_in_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --niosII_openMac_clock_1_in_beginbursttransfer_internal begin burst transfer, which is an e_assign
  niosII_openMac_clock_1_in_beginbursttransfer_internal <= niosII_openMac_clock_1_in_begins_xfer;
  --niosII_openMac_clock_1_in_read assignment, which is an e_mux
  niosII_openMac_clock_1_in_read <= internal_pcp_cpu_data_master_granted_niosII_openMac_clock_1_in AND pcp_cpu_data_master_read;
  --niosII_openMac_clock_1_in_write assignment, which is an e_mux
  niosII_openMac_clock_1_in_write <= internal_pcp_cpu_data_master_granted_niosII_openMac_clock_1_in AND pcp_cpu_data_master_write;
  --niosII_openMac_clock_1_in_address mux, which is an e_mux
  niosII_openMac_clock_1_in_address <= pcp_cpu_data_master_address_to_slave (2 DOWNTO 0);
  --slaveid niosII_openMac_clock_1_in_nativeaddress nativeaddress mux, which is an e_mux
  niosII_openMac_clock_1_in_nativeaddress <= Vector_To_Std_Logic(A_SRL(pcp_cpu_data_master_address_to_slave,std_logic_vector'("00000000000000000000000000000010")));
  --d1_niosII_openMac_clock_1_in_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_niosII_openMac_clock_1_in_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_niosII_openMac_clock_1_in_end_xfer <= niosII_openMac_clock_1_in_end_xfer;
    end if;

  end process;

  --niosII_openMac_clock_1_in_waits_for_read in a cycle, which is an e_mux
  niosII_openMac_clock_1_in_waits_for_read <= niosII_openMac_clock_1_in_in_a_read_cycle AND internal_niosII_openMac_clock_1_in_waitrequest_from_sa;
  --niosII_openMac_clock_1_in_in_a_read_cycle assignment, which is an e_assign
  niosII_openMac_clock_1_in_in_a_read_cycle <= internal_pcp_cpu_data_master_granted_niosII_openMac_clock_1_in AND pcp_cpu_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= niosII_openMac_clock_1_in_in_a_read_cycle;
  --niosII_openMac_clock_1_in_waits_for_write in a cycle, which is an e_mux
  niosII_openMac_clock_1_in_waits_for_write <= niosII_openMac_clock_1_in_in_a_write_cycle AND internal_niosII_openMac_clock_1_in_waitrequest_from_sa;
  --niosII_openMac_clock_1_in_in_a_write_cycle assignment, which is an e_assign
  niosII_openMac_clock_1_in_in_a_write_cycle <= internal_pcp_cpu_data_master_granted_niosII_openMac_clock_1_in AND pcp_cpu_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= niosII_openMac_clock_1_in_in_a_write_cycle;
  wait_for_niosII_openMac_clock_1_in_counter <= std_logic'('0');
  --niosII_openMac_clock_1_in_byteenable byte enable port mux, which is an e_mux
  niosII_openMac_clock_1_in_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_pcp_cpu_data_master_granted_niosII_openMac_clock_1_in)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (pcp_cpu_data_master_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))), 4);
  --vhdl renameroo for output signals
  niosII_openMac_clock_1_in_waitrequest_from_sa <= internal_niosII_openMac_clock_1_in_waitrequest_from_sa;
  --vhdl renameroo for output signals
  pcp_cpu_data_master_granted_niosII_openMac_clock_1_in <= internal_pcp_cpu_data_master_granted_niosII_openMac_clock_1_in;
  --vhdl renameroo for output signals
  pcp_cpu_data_master_qualified_request_niosII_openMac_clock_1_in <= internal_pcp_cpu_data_master_qualified_request_niosII_openMac_clock_1_in;
  --vhdl renameroo for output signals
  pcp_cpu_data_master_requests_niosII_openMac_clock_1_in <= internal_pcp_cpu_data_master_requests_niosII_openMac_clock_1_in;
--synthesis translate_off
    --niosII_openMac_clock_1/in enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity niosII_openMac_clock_1_out_arbitrator is 
        port (
              -- inputs:
                 signal OpenMAC_0_CMP_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal clk : IN STD_LOGIC;
                 signal d1_OpenMAC_0_CMP_end_xfer : IN STD_LOGIC;
                 signal niosII_openMac_clock_1_out_address : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal niosII_openMac_clock_1_out_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal niosII_openMac_clock_1_out_granted_OpenMAC_0_CMP : IN STD_LOGIC;
                 signal niosII_openMac_clock_1_out_qualified_request_OpenMAC_0_CMP : IN STD_LOGIC;
                 signal niosII_openMac_clock_1_out_read : IN STD_LOGIC;
                 signal niosII_openMac_clock_1_out_read_data_valid_OpenMAC_0_CMP : IN STD_LOGIC;
                 signal niosII_openMac_clock_1_out_requests_OpenMAC_0_CMP : IN STD_LOGIC;
                 signal niosII_openMac_clock_1_out_write : IN STD_LOGIC;
                 signal niosII_openMac_clock_1_out_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal niosII_openMac_clock_1_out_address_to_slave : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal niosII_openMac_clock_1_out_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal niosII_openMac_clock_1_out_reset_n : OUT STD_LOGIC;
                 signal niosII_openMac_clock_1_out_waitrequest : OUT STD_LOGIC
              );
end entity niosII_openMac_clock_1_out_arbitrator;


architecture europa of niosII_openMac_clock_1_out_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal internal_niosII_openMac_clock_1_out_address_to_slave :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal internal_niosII_openMac_clock_1_out_waitrequest :  STD_LOGIC;
                signal niosII_openMac_clock_1_out_address_last_time :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal niosII_openMac_clock_1_out_byteenable_last_time :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_openMac_clock_1_out_read_last_time :  STD_LOGIC;
                signal niosII_openMac_clock_1_out_run :  STD_LOGIC;
                signal niosII_openMac_clock_1_out_write_last_time :  STD_LOGIC;
                signal niosII_openMac_clock_1_out_writedata_last_time :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal r_0 :  STD_LOGIC;

begin

  --r_0 master_run cascaded wait assignment, which is an e_assign
  r_0 <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000001") AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT niosII_openMac_clock_1_out_qualified_request_OpenMAC_0_CMP OR NOT niosII_openMac_clock_1_out_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT d1_OpenMAC_0_CMP_end_xfer)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(niosII_openMac_clock_1_out_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT niosII_openMac_clock_1_out_qualified_request_OpenMAC_0_CMP OR NOT niosII_openMac_clock_1_out_write)))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(niosII_openMac_clock_1_out_write)))))))));
  --cascaded wait assignment, which is an e_assign
  niosII_openMac_clock_1_out_run <= r_0;
  --optimize select-logic by passing only those address bits which matter.
  internal_niosII_openMac_clock_1_out_address_to_slave <= niosII_openMac_clock_1_out_address;
  --niosII_openMac_clock_1/out readdata mux, which is an e_mux
  niosII_openMac_clock_1_out_readdata <= OpenMAC_0_CMP_readdata_from_sa;
  --actual waitrequest port, which is an e_assign
  internal_niosII_openMac_clock_1_out_waitrequest <= NOT niosII_openMac_clock_1_out_run;
  --niosII_openMac_clock_1_out_reset_n assignment, which is an e_assign
  niosII_openMac_clock_1_out_reset_n <= reset_n;
  --vhdl renameroo for output signals
  niosII_openMac_clock_1_out_address_to_slave <= internal_niosII_openMac_clock_1_out_address_to_slave;
  --vhdl renameroo for output signals
  niosII_openMac_clock_1_out_waitrequest <= internal_niosII_openMac_clock_1_out_waitrequest;
--synthesis translate_off
    --niosII_openMac_clock_1_out_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_openMac_clock_1_out_address_last_time <= std_logic_vector'("000");
      elsif clk'event and clk = '1' then
        niosII_openMac_clock_1_out_address_last_time <= niosII_openMac_clock_1_out_address;
      end if;

    end process;

    --niosII_openMac_clock_1/out waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_niosII_openMac_clock_1_out_waitrequest AND ((niosII_openMac_clock_1_out_read OR niosII_openMac_clock_1_out_write));
      end if;

    end process;

    --niosII_openMac_clock_1_out_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line21 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((niosII_openMac_clock_1_out_address /= niosII_openMac_clock_1_out_address_last_time))))) = '1' then 
          write(write_line21, now);
          write(write_line21, string'(": "));
          write(write_line21, string'("niosII_openMac_clock_1_out_address did not heed wait!!!"));
          write(output, write_line21.all);
          deallocate (write_line21);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_openMac_clock_1_out_byteenable check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_openMac_clock_1_out_byteenable_last_time <= std_logic_vector'("0000");
      elsif clk'event and clk = '1' then
        niosII_openMac_clock_1_out_byteenable_last_time <= niosII_openMac_clock_1_out_byteenable;
      end if;

    end process;

    --niosII_openMac_clock_1_out_byteenable matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line22 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((niosII_openMac_clock_1_out_byteenable /= niosII_openMac_clock_1_out_byteenable_last_time))))) = '1' then 
          write(write_line22, now);
          write(write_line22, string'(": "));
          write(write_line22, string'("niosII_openMac_clock_1_out_byteenable did not heed wait!!!"));
          write(output, write_line22.all);
          deallocate (write_line22);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_openMac_clock_1_out_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_openMac_clock_1_out_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        niosII_openMac_clock_1_out_read_last_time <= niosII_openMac_clock_1_out_read;
      end if;

    end process;

    --niosII_openMac_clock_1_out_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line23 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(niosII_openMac_clock_1_out_read) /= std_logic'(niosII_openMac_clock_1_out_read_last_time)))))) = '1' then 
          write(write_line23, now);
          write(write_line23, string'(": "));
          write(write_line23, string'("niosII_openMac_clock_1_out_read did not heed wait!!!"));
          write(output, write_line23.all);
          deallocate (write_line23);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_openMac_clock_1_out_write check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_openMac_clock_1_out_write_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        niosII_openMac_clock_1_out_write_last_time <= niosII_openMac_clock_1_out_write;
      end if;

    end process;

    --niosII_openMac_clock_1_out_write matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line24 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(niosII_openMac_clock_1_out_write) /= std_logic'(niosII_openMac_clock_1_out_write_last_time)))))) = '1' then 
          write(write_line24, now);
          write(write_line24, string'(": "));
          write(write_line24, string'("niosII_openMac_clock_1_out_write did not heed wait!!!"));
          write(output, write_line24.all);
          deallocate (write_line24);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_openMac_clock_1_out_writedata check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_openMac_clock_1_out_writedata_last_time <= std_logic_vector'("00000000000000000000000000000000");
      elsif clk'event and clk = '1' then
        niosII_openMac_clock_1_out_writedata_last_time <= niosII_openMac_clock_1_out_writedata;
      end if;

    end process;

    --niosII_openMac_clock_1_out_writedata matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line25 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((active_and_waiting_last_time AND to_std_logic(((niosII_openMac_clock_1_out_writedata /= niosII_openMac_clock_1_out_writedata_last_time)))) AND niosII_openMac_clock_1_out_write)) = '1' then 
          write(write_line25, now);
          write(write_line25, string'(": "));
          write(write_line25, string'("niosII_openMac_clock_1_out_writedata did not heed wait!!!"));
          write(output, write_line25.all);
          deallocate (write_line25);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity niosII_openMac_clock_2_in_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal niosII_openMac_clock_2_in_endofpacket : IN STD_LOGIC;
                 signal niosII_openMac_clock_2_in_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal niosII_openMac_clock_2_in_waitrequest : IN STD_LOGIC;
                 signal pcp_cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (25 DOWNTO 0);
                 signal pcp_cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal pcp_cpu_data_master_dbs_address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal pcp_cpu_data_master_dbs_write_16 : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal pcp_cpu_data_master_no_byte_enables_and_last_term : IN STD_LOGIC;
                 signal pcp_cpu_data_master_read : IN STD_LOGIC;
                 signal pcp_cpu_data_master_waitrequest : IN STD_LOGIC;
                 signal pcp_cpu_data_master_write : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal d1_niosII_openMac_clock_2_in_end_xfer : OUT STD_LOGIC;
                 signal niosII_openMac_clock_2_in_address : OUT STD_LOGIC_VECTOR (12 DOWNTO 0);
                 signal niosII_openMac_clock_2_in_byteenable : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal niosII_openMac_clock_2_in_endofpacket_from_sa : OUT STD_LOGIC;
                 signal niosII_openMac_clock_2_in_nativeaddress : OUT STD_LOGIC_VECTOR (11 DOWNTO 0);
                 signal niosII_openMac_clock_2_in_read : OUT STD_LOGIC;
                 signal niosII_openMac_clock_2_in_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal niosII_openMac_clock_2_in_reset_n : OUT STD_LOGIC;
                 signal niosII_openMac_clock_2_in_waitrequest_from_sa : OUT STD_LOGIC;
                 signal niosII_openMac_clock_2_in_write : OUT STD_LOGIC;
                 signal niosII_openMac_clock_2_in_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal pcp_cpu_data_master_byteenable_niosII_openMac_clock_2_in : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal pcp_cpu_data_master_granted_niosII_openMac_clock_2_in : OUT STD_LOGIC;
                 signal pcp_cpu_data_master_qualified_request_niosII_openMac_clock_2_in : OUT STD_LOGIC;
                 signal pcp_cpu_data_master_read_data_valid_niosII_openMac_clock_2_in : OUT STD_LOGIC;
                 signal pcp_cpu_data_master_requests_niosII_openMac_clock_2_in : OUT STD_LOGIC
              );
end entity niosII_openMac_clock_2_in_arbitrator;


architecture europa of niosII_openMac_clock_2_in_arbitrator is
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_niosII_openMac_clock_2_in :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_niosII_openMac_clock_2_in_waitrequest_from_sa :  STD_LOGIC;
                signal internal_pcp_cpu_data_master_byteenable_niosII_openMac_clock_2_in :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal internal_pcp_cpu_data_master_granted_niosII_openMac_clock_2_in :  STD_LOGIC;
                signal internal_pcp_cpu_data_master_qualified_request_niosII_openMac_clock_2_in :  STD_LOGIC;
                signal internal_pcp_cpu_data_master_requests_niosII_openMac_clock_2_in :  STD_LOGIC;
                signal niosII_openMac_clock_2_in_allgrants :  STD_LOGIC;
                signal niosII_openMac_clock_2_in_allow_new_arb_cycle :  STD_LOGIC;
                signal niosII_openMac_clock_2_in_any_bursting_master_saved_grant :  STD_LOGIC;
                signal niosII_openMac_clock_2_in_any_continuerequest :  STD_LOGIC;
                signal niosII_openMac_clock_2_in_arb_counter_enable :  STD_LOGIC;
                signal niosII_openMac_clock_2_in_arb_share_counter :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal niosII_openMac_clock_2_in_arb_share_counter_next_value :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal niosII_openMac_clock_2_in_arb_share_set_values :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal niosII_openMac_clock_2_in_beginbursttransfer_internal :  STD_LOGIC;
                signal niosII_openMac_clock_2_in_begins_xfer :  STD_LOGIC;
                signal niosII_openMac_clock_2_in_end_xfer :  STD_LOGIC;
                signal niosII_openMac_clock_2_in_firsttransfer :  STD_LOGIC;
                signal niosII_openMac_clock_2_in_grant_vector :  STD_LOGIC;
                signal niosII_openMac_clock_2_in_in_a_read_cycle :  STD_LOGIC;
                signal niosII_openMac_clock_2_in_in_a_write_cycle :  STD_LOGIC;
                signal niosII_openMac_clock_2_in_master_qreq_vector :  STD_LOGIC;
                signal niosII_openMac_clock_2_in_non_bursting_master_requests :  STD_LOGIC;
                signal niosII_openMac_clock_2_in_reg_firsttransfer :  STD_LOGIC;
                signal niosII_openMac_clock_2_in_slavearbiterlockenable :  STD_LOGIC;
                signal niosII_openMac_clock_2_in_slavearbiterlockenable2 :  STD_LOGIC;
                signal niosII_openMac_clock_2_in_unreg_firsttransfer :  STD_LOGIC;
                signal niosII_openMac_clock_2_in_waits_for_read :  STD_LOGIC;
                signal niosII_openMac_clock_2_in_waits_for_write :  STD_LOGIC;
                signal pcp_cpu_data_master_arbiterlock :  STD_LOGIC;
                signal pcp_cpu_data_master_arbiterlock2 :  STD_LOGIC;
                signal pcp_cpu_data_master_byteenable_niosII_openMac_clock_2_in_segment_0 :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal pcp_cpu_data_master_byteenable_niosII_openMac_clock_2_in_segment_1 :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal pcp_cpu_data_master_continuerequest :  STD_LOGIC;
                signal pcp_cpu_data_master_saved_grant_niosII_openMac_clock_2_in :  STD_LOGIC;
                signal wait_for_niosII_openMac_clock_2_in_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT niosII_openMac_clock_2_in_end_xfer;
    end if;

  end process;

  niosII_openMac_clock_2_in_begins_xfer <= NOT d1_reasons_to_wait AND (internal_pcp_cpu_data_master_qualified_request_niosII_openMac_clock_2_in);
  --assign niosII_openMac_clock_2_in_readdata_from_sa = niosII_openMac_clock_2_in_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  niosII_openMac_clock_2_in_readdata_from_sa <= niosII_openMac_clock_2_in_readdata;
  internal_pcp_cpu_data_master_requests_niosII_openMac_clock_2_in <= to_std_logic(((Std_Logic_Vector'(pcp_cpu_data_master_address_to_slave(25 DOWNTO 13) & std_logic_vector'("0000000000000")) = std_logic_vector'("00000000000010000000000000")))) AND ((pcp_cpu_data_master_read OR pcp_cpu_data_master_write));
  --assign niosII_openMac_clock_2_in_waitrequest_from_sa = niosII_openMac_clock_2_in_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_niosII_openMac_clock_2_in_waitrequest_from_sa <= niosII_openMac_clock_2_in_waitrequest;
  --niosII_openMac_clock_2_in_arb_share_counter set values, which is an e_mux
  niosII_openMac_clock_2_in_arb_share_set_values <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_pcp_cpu_data_master_granted_niosII_openMac_clock_2_in)) = '1'), std_logic_vector'("00000000000000000000000000000010"), std_logic_vector'("00000000000000000000000000000001")), 2);
  --niosII_openMac_clock_2_in_non_bursting_master_requests mux, which is an e_mux
  niosII_openMac_clock_2_in_non_bursting_master_requests <= internal_pcp_cpu_data_master_requests_niosII_openMac_clock_2_in;
  --niosII_openMac_clock_2_in_any_bursting_master_saved_grant mux, which is an e_mux
  niosII_openMac_clock_2_in_any_bursting_master_saved_grant <= std_logic'('0');
  --niosII_openMac_clock_2_in_arb_share_counter_next_value assignment, which is an e_assign
  niosII_openMac_clock_2_in_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(niosII_openMac_clock_2_in_firsttransfer) = '1'), (((std_logic_vector'("0000000000000000000000000000000") & (niosII_openMac_clock_2_in_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(niosII_openMac_clock_2_in_arb_share_counter)) = '1'), (((std_logic_vector'("0000000000000000000000000000000") & (niosII_openMac_clock_2_in_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 2);
  --niosII_openMac_clock_2_in_allgrants all slave grants, which is an e_mux
  niosII_openMac_clock_2_in_allgrants <= niosII_openMac_clock_2_in_grant_vector;
  --niosII_openMac_clock_2_in_end_xfer assignment, which is an e_assign
  niosII_openMac_clock_2_in_end_xfer <= NOT ((niosII_openMac_clock_2_in_waits_for_read OR niosII_openMac_clock_2_in_waits_for_write));
  --end_xfer_arb_share_counter_term_niosII_openMac_clock_2_in arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_niosII_openMac_clock_2_in <= niosII_openMac_clock_2_in_end_xfer AND (((NOT niosII_openMac_clock_2_in_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --niosII_openMac_clock_2_in_arb_share_counter arbitration counter enable, which is an e_assign
  niosII_openMac_clock_2_in_arb_counter_enable <= ((end_xfer_arb_share_counter_term_niosII_openMac_clock_2_in AND niosII_openMac_clock_2_in_allgrants)) OR ((end_xfer_arb_share_counter_term_niosII_openMac_clock_2_in AND NOT niosII_openMac_clock_2_in_non_bursting_master_requests));
  --niosII_openMac_clock_2_in_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_openMac_clock_2_in_arb_share_counter <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      if std_logic'(niosII_openMac_clock_2_in_arb_counter_enable) = '1' then 
        niosII_openMac_clock_2_in_arb_share_counter <= niosII_openMac_clock_2_in_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --niosII_openMac_clock_2_in_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_openMac_clock_2_in_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((niosII_openMac_clock_2_in_master_qreq_vector AND end_xfer_arb_share_counter_term_niosII_openMac_clock_2_in)) OR ((end_xfer_arb_share_counter_term_niosII_openMac_clock_2_in AND NOT niosII_openMac_clock_2_in_non_bursting_master_requests)))) = '1' then 
        niosII_openMac_clock_2_in_slavearbiterlockenable <= or_reduce(niosII_openMac_clock_2_in_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --pcp_cpu/data_master niosII_openMac_clock_2/in arbiterlock, which is an e_assign
  pcp_cpu_data_master_arbiterlock <= niosII_openMac_clock_2_in_slavearbiterlockenable AND pcp_cpu_data_master_continuerequest;
  --niosII_openMac_clock_2_in_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  niosII_openMac_clock_2_in_slavearbiterlockenable2 <= or_reduce(niosII_openMac_clock_2_in_arb_share_counter_next_value);
  --pcp_cpu/data_master niosII_openMac_clock_2/in arbiterlock2, which is an e_assign
  pcp_cpu_data_master_arbiterlock2 <= niosII_openMac_clock_2_in_slavearbiterlockenable2 AND pcp_cpu_data_master_continuerequest;
  --niosII_openMac_clock_2_in_any_continuerequest at least one master continues requesting, which is an e_assign
  niosII_openMac_clock_2_in_any_continuerequest <= std_logic'('1');
  --pcp_cpu_data_master_continuerequest continued request, which is an e_assign
  pcp_cpu_data_master_continuerequest <= std_logic'('1');
  internal_pcp_cpu_data_master_qualified_request_niosII_openMac_clock_2_in <= internal_pcp_cpu_data_master_requests_niosII_openMac_clock_2_in AND NOT ((((pcp_cpu_data_master_read AND (NOT pcp_cpu_data_master_waitrequest))) OR (((((NOT pcp_cpu_data_master_waitrequest OR pcp_cpu_data_master_no_byte_enables_and_last_term) OR NOT(or_reduce(internal_pcp_cpu_data_master_byteenable_niosII_openMac_clock_2_in)))) AND pcp_cpu_data_master_write))));
  --niosII_openMac_clock_2_in_writedata mux, which is an e_mux
  niosII_openMac_clock_2_in_writedata <= pcp_cpu_data_master_dbs_write_16;
  --assign niosII_openMac_clock_2_in_endofpacket_from_sa = niosII_openMac_clock_2_in_endofpacket so that symbol knows where to group signals which may go to master only, which is an e_assign
  niosII_openMac_clock_2_in_endofpacket_from_sa <= niosII_openMac_clock_2_in_endofpacket;
  --master is always granted when requested
  internal_pcp_cpu_data_master_granted_niosII_openMac_clock_2_in <= internal_pcp_cpu_data_master_qualified_request_niosII_openMac_clock_2_in;
  --pcp_cpu/data_master saved-grant niosII_openMac_clock_2/in, which is an e_assign
  pcp_cpu_data_master_saved_grant_niosII_openMac_clock_2_in <= internal_pcp_cpu_data_master_requests_niosII_openMac_clock_2_in;
  --allow new arb cycle for niosII_openMac_clock_2/in, which is an e_assign
  niosII_openMac_clock_2_in_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  niosII_openMac_clock_2_in_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  niosII_openMac_clock_2_in_master_qreq_vector <= std_logic'('1');
  --niosII_openMac_clock_2_in_reset_n assignment, which is an e_assign
  niosII_openMac_clock_2_in_reset_n <= reset_n;
  --niosII_openMac_clock_2_in_firsttransfer first transaction, which is an e_assign
  niosII_openMac_clock_2_in_firsttransfer <= A_WE_StdLogic((std_logic'(niosII_openMac_clock_2_in_begins_xfer) = '1'), niosII_openMac_clock_2_in_unreg_firsttransfer, niosII_openMac_clock_2_in_reg_firsttransfer);
  --niosII_openMac_clock_2_in_unreg_firsttransfer first transaction, which is an e_assign
  niosII_openMac_clock_2_in_unreg_firsttransfer <= NOT ((niosII_openMac_clock_2_in_slavearbiterlockenable AND niosII_openMac_clock_2_in_any_continuerequest));
  --niosII_openMac_clock_2_in_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_openMac_clock_2_in_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(niosII_openMac_clock_2_in_begins_xfer) = '1' then 
        niosII_openMac_clock_2_in_reg_firsttransfer <= niosII_openMac_clock_2_in_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --niosII_openMac_clock_2_in_beginbursttransfer_internal begin burst transfer, which is an e_assign
  niosII_openMac_clock_2_in_beginbursttransfer_internal <= niosII_openMac_clock_2_in_begins_xfer;
  --niosII_openMac_clock_2_in_read assignment, which is an e_mux
  niosII_openMac_clock_2_in_read <= internal_pcp_cpu_data_master_granted_niosII_openMac_clock_2_in AND pcp_cpu_data_master_read;
  --niosII_openMac_clock_2_in_write assignment, which is an e_mux
  niosII_openMac_clock_2_in_write <= internal_pcp_cpu_data_master_granted_niosII_openMac_clock_2_in AND pcp_cpu_data_master_write;
  --niosII_openMac_clock_2_in_address mux, which is an e_mux
  niosII_openMac_clock_2_in_address <= A_EXT (Std_Logic_Vector'(A_SRL(pcp_cpu_data_master_address_to_slave,std_logic_vector'("00000000000000000000000000000010")) & A_ToStdLogicVector(pcp_cpu_data_master_dbs_address(1)) & A_ToStdLogicVector(std_logic'('0'))), 13);
  --slaveid niosII_openMac_clock_2_in_nativeaddress nativeaddress mux, which is an e_mux
  niosII_openMac_clock_2_in_nativeaddress <= A_EXT (A_SRL(pcp_cpu_data_master_address_to_slave,std_logic_vector'("00000000000000000000000000000010")), 12);
  --d1_niosII_openMac_clock_2_in_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_niosII_openMac_clock_2_in_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_niosII_openMac_clock_2_in_end_xfer <= niosII_openMac_clock_2_in_end_xfer;
    end if;

  end process;

  --niosII_openMac_clock_2_in_waits_for_read in a cycle, which is an e_mux
  niosII_openMac_clock_2_in_waits_for_read <= niosII_openMac_clock_2_in_in_a_read_cycle AND internal_niosII_openMac_clock_2_in_waitrequest_from_sa;
  --niosII_openMac_clock_2_in_in_a_read_cycle assignment, which is an e_assign
  niosII_openMac_clock_2_in_in_a_read_cycle <= internal_pcp_cpu_data_master_granted_niosII_openMac_clock_2_in AND pcp_cpu_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= niosII_openMac_clock_2_in_in_a_read_cycle;
  --niosII_openMac_clock_2_in_waits_for_write in a cycle, which is an e_mux
  niosII_openMac_clock_2_in_waits_for_write <= niosII_openMac_clock_2_in_in_a_write_cycle AND internal_niosII_openMac_clock_2_in_waitrequest_from_sa;
  --niosII_openMac_clock_2_in_in_a_write_cycle assignment, which is an e_assign
  niosII_openMac_clock_2_in_in_a_write_cycle <= internal_pcp_cpu_data_master_granted_niosII_openMac_clock_2_in AND pcp_cpu_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= niosII_openMac_clock_2_in_in_a_write_cycle;
  wait_for_niosII_openMac_clock_2_in_counter <= std_logic'('0');
  --niosII_openMac_clock_2_in_byteenable byte enable port mux, which is an e_mux
  niosII_openMac_clock_2_in_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_pcp_cpu_data_master_granted_niosII_openMac_clock_2_in)) = '1'), (std_logic_vector'("000000000000000000000000000000") & (internal_pcp_cpu_data_master_byteenable_niosII_openMac_clock_2_in)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))), 2);
  (pcp_cpu_data_master_byteenable_niosII_openMac_clock_2_in_segment_1(1), pcp_cpu_data_master_byteenable_niosII_openMac_clock_2_in_segment_1(0), pcp_cpu_data_master_byteenable_niosII_openMac_clock_2_in_segment_0(1), pcp_cpu_data_master_byteenable_niosII_openMac_clock_2_in_segment_0(0)) <= pcp_cpu_data_master_byteenable;
  internal_pcp_cpu_data_master_byteenable_niosII_openMac_clock_2_in <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pcp_cpu_data_master_dbs_address(1)))) = std_logic_vector'("00000000000000000000000000000000"))), pcp_cpu_data_master_byteenable_niosII_openMac_clock_2_in_segment_0, pcp_cpu_data_master_byteenable_niosII_openMac_clock_2_in_segment_1);
  --vhdl renameroo for output signals
  niosII_openMac_clock_2_in_waitrequest_from_sa <= internal_niosII_openMac_clock_2_in_waitrequest_from_sa;
  --vhdl renameroo for output signals
  pcp_cpu_data_master_byteenable_niosII_openMac_clock_2_in <= internal_pcp_cpu_data_master_byteenable_niosII_openMac_clock_2_in;
  --vhdl renameroo for output signals
  pcp_cpu_data_master_granted_niosII_openMac_clock_2_in <= internal_pcp_cpu_data_master_granted_niosII_openMac_clock_2_in;
  --vhdl renameroo for output signals
  pcp_cpu_data_master_qualified_request_niosII_openMac_clock_2_in <= internal_pcp_cpu_data_master_qualified_request_niosII_openMac_clock_2_in;
  --vhdl renameroo for output signals
  pcp_cpu_data_master_requests_niosII_openMac_clock_2_in <= internal_pcp_cpu_data_master_requests_niosII_openMac_clock_2_in;
--synthesis translate_off
    --niosII_openMac_clock_2/in enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity niosII_openMac_clock_2_out_arbitrator is 
        port (
              -- inputs:
                 signal OpenMAC_0_REG_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal clk : IN STD_LOGIC;
                 signal d1_OpenMAC_0_REG_end_xfer : IN STD_LOGIC;
                 signal niosII_openMac_clock_2_out_address : IN STD_LOGIC_VECTOR (12 DOWNTO 0);
                 signal niosII_openMac_clock_2_out_byteenable : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal niosII_openMac_clock_2_out_granted_OpenMAC_0_REG : IN STD_LOGIC;
                 signal niosII_openMac_clock_2_out_qualified_request_OpenMAC_0_REG : IN STD_LOGIC;
                 signal niosII_openMac_clock_2_out_read : IN STD_LOGIC;
                 signal niosII_openMac_clock_2_out_read_data_valid_OpenMAC_0_REG : IN STD_LOGIC;
                 signal niosII_openMac_clock_2_out_requests_OpenMAC_0_REG : IN STD_LOGIC;
                 signal niosII_openMac_clock_2_out_write : IN STD_LOGIC;
                 signal niosII_openMac_clock_2_out_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal niosII_openMac_clock_2_out_address_to_slave : OUT STD_LOGIC_VECTOR (12 DOWNTO 0);
                 signal niosII_openMac_clock_2_out_readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal niosII_openMac_clock_2_out_reset_n : OUT STD_LOGIC;
                 signal niosII_openMac_clock_2_out_waitrequest : OUT STD_LOGIC
              );
end entity niosII_openMac_clock_2_out_arbitrator;


architecture europa of niosII_openMac_clock_2_out_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal internal_niosII_openMac_clock_2_out_address_to_slave :  STD_LOGIC_VECTOR (12 DOWNTO 0);
                signal internal_niosII_openMac_clock_2_out_waitrequest :  STD_LOGIC;
                signal niosII_openMac_clock_2_out_address_last_time :  STD_LOGIC_VECTOR (12 DOWNTO 0);
                signal niosII_openMac_clock_2_out_byteenable_last_time :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal niosII_openMac_clock_2_out_read_last_time :  STD_LOGIC;
                signal niosII_openMac_clock_2_out_run :  STD_LOGIC;
                signal niosII_openMac_clock_2_out_write_last_time :  STD_LOGIC;
                signal niosII_openMac_clock_2_out_writedata_last_time :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal r_0 :  STD_LOGIC;

begin

  --r_0 master_run cascaded wait assignment, which is an e_assign
  r_0 <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000001") AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT niosII_openMac_clock_2_out_qualified_request_OpenMAC_0_REG OR NOT niosII_openMac_clock_2_out_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT d1_OpenMAC_0_REG_end_xfer)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(niosII_openMac_clock_2_out_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT niosII_openMac_clock_2_out_qualified_request_OpenMAC_0_REG OR NOT niosII_openMac_clock_2_out_write)))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(niosII_openMac_clock_2_out_write)))))))));
  --cascaded wait assignment, which is an e_assign
  niosII_openMac_clock_2_out_run <= r_0;
  --optimize select-logic by passing only those address bits which matter.
  internal_niosII_openMac_clock_2_out_address_to_slave <= niosII_openMac_clock_2_out_address;
  --niosII_openMac_clock_2/out readdata mux, which is an e_mux
  niosII_openMac_clock_2_out_readdata <= OpenMAC_0_REG_readdata_from_sa;
  --actual waitrequest port, which is an e_assign
  internal_niosII_openMac_clock_2_out_waitrequest <= NOT niosII_openMac_clock_2_out_run;
  --niosII_openMac_clock_2_out_reset_n assignment, which is an e_assign
  niosII_openMac_clock_2_out_reset_n <= reset_n;
  --vhdl renameroo for output signals
  niosII_openMac_clock_2_out_address_to_slave <= internal_niosII_openMac_clock_2_out_address_to_slave;
  --vhdl renameroo for output signals
  niosII_openMac_clock_2_out_waitrequest <= internal_niosII_openMac_clock_2_out_waitrequest;
--synthesis translate_off
    --niosII_openMac_clock_2_out_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_openMac_clock_2_out_address_last_time <= std_logic_vector'("0000000000000");
      elsif clk'event and clk = '1' then
        niosII_openMac_clock_2_out_address_last_time <= niosII_openMac_clock_2_out_address;
      end if;

    end process;

    --niosII_openMac_clock_2/out waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_niosII_openMac_clock_2_out_waitrequest AND ((niosII_openMac_clock_2_out_read OR niosII_openMac_clock_2_out_write));
      end if;

    end process;

    --niosII_openMac_clock_2_out_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line26 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((niosII_openMac_clock_2_out_address /= niosII_openMac_clock_2_out_address_last_time))))) = '1' then 
          write(write_line26, now);
          write(write_line26, string'(": "));
          write(write_line26, string'("niosII_openMac_clock_2_out_address did not heed wait!!!"));
          write(output, write_line26.all);
          deallocate (write_line26);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_openMac_clock_2_out_byteenable check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_openMac_clock_2_out_byteenable_last_time <= std_logic_vector'("00");
      elsif clk'event and clk = '1' then
        niosII_openMac_clock_2_out_byteenable_last_time <= niosII_openMac_clock_2_out_byteenable;
      end if;

    end process;

    --niosII_openMac_clock_2_out_byteenable matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line27 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((niosII_openMac_clock_2_out_byteenable /= niosII_openMac_clock_2_out_byteenable_last_time))))) = '1' then 
          write(write_line27, now);
          write(write_line27, string'(": "));
          write(write_line27, string'("niosII_openMac_clock_2_out_byteenable did not heed wait!!!"));
          write(output, write_line27.all);
          deallocate (write_line27);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_openMac_clock_2_out_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_openMac_clock_2_out_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        niosII_openMac_clock_2_out_read_last_time <= niosII_openMac_clock_2_out_read;
      end if;

    end process;

    --niosII_openMac_clock_2_out_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line28 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(niosII_openMac_clock_2_out_read) /= std_logic'(niosII_openMac_clock_2_out_read_last_time)))))) = '1' then 
          write(write_line28, now);
          write(write_line28, string'(": "));
          write(write_line28, string'("niosII_openMac_clock_2_out_read did not heed wait!!!"));
          write(output, write_line28.all);
          deallocate (write_line28);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_openMac_clock_2_out_write check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_openMac_clock_2_out_write_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        niosII_openMac_clock_2_out_write_last_time <= niosII_openMac_clock_2_out_write;
      end if;

    end process;

    --niosII_openMac_clock_2_out_write matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line29 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(niosII_openMac_clock_2_out_write) /= std_logic'(niosII_openMac_clock_2_out_write_last_time)))))) = '1' then 
          write(write_line29, now);
          write(write_line29, string'(": "));
          write(write_line29, string'("niosII_openMac_clock_2_out_write did not heed wait!!!"));
          write(output, write_line29.all);
          deallocate (write_line29);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_openMac_clock_2_out_writedata check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_openMac_clock_2_out_writedata_last_time <= std_logic_vector'("0000000000000000");
      elsif clk'event and clk = '1' then
        niosII_openMac_clock_2_out_writedata_last_time <= niosII_openMac_clock_2_out_writedata;
      end if;

    end process;

    --niosII_openMac_clock_2_out_writedata matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line30 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((active_and_waiting_last_time AND to_std_logic(((niosII_openMac_clock_2_out_writedata /= niosII_openMac_clock_2_out_writedata_last_time)))) AND niosII_openMac_clock_2_out_write)) = '1' then 
          write(write_line30, now);
          write(write_line30, string'(": "));
          write(write_line30, string'("niosII_openMac_clock_2_out_writedata did not heed wait!!!"));
          write(output, write_line30.all);
          deallocate (write_line30);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity niosII_openMac_clock_3_in_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal niosII_openMac_clock_3_in_endofpacket : IN STD_LOGIC;
                 signal niosII_openMac_clock_3_in_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal niosII_openMac_clock_3_in_waitrequest : IN STD_LOGIC;
                 signal pcp_cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (25 DOWNTO 0);
                 signal pcp_cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal pcp_cpu_data_master_read : IN STD_LOGIC;
                 signal pcp_cpu_data_master_waitrequest : IN STD_LOGIC;
                 signal pcp_cpu_data_master_write : IN STD_LOGIC;
                 signal pcp_cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal d1_niosII_openMac_clock_3_in_end_xfer : OUT STD_LOGIC;
                 signal niosII_openMac_clock_3_in_address : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal niosII_openMac_clock_3_in_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal niosII_openMac_clock_3_in_endofpacket_from_sa : OUT STD_LOGIC;
                 signal niosII_openMac_clock_3_in_nativeaddress : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal niosII_openMac_clock_3_in_read : OUT STD_LOGIC;
                 signal niosII_openMac_clock_3_in_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal niosII_openMac_clock_3_in_reset_n : OUT STD_LOGIC;
                 signal niosII_openMac_clock_3_in_waitrequest_from_sa : OUT STD_LOGIC;
                 signal niosII_openMac_clock_3_in_write : OUT STD_LOGIC;
                 signal niosII_openMac_clock_3_in_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal pcp_cpu_data_master_granted_niosII_openMac_clock_3_in : OUT STD_LOGIC;
                 signal pcp_cpu_data_master_qualified_request_niosII_openMac_clock_3_in : OUT STD_LOGIC;
                 signal pcp_cpu_data_master_read_data_valid_niosII_openMac_clock_3_in : OUT STD_LOGIC;
                 signal pcp_cpu_data_master_requests_niosII_openMac_clock_3_in : OUT STD_LOGIC
              );
end entity niosII_openMac_clock_3_in_arbitrator;


architecture europa of niosII_openMac_clock_3_in_arbitrator is
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_niosII_openMac_clock_3_in :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_niosII_openMac_clock_3_in_waitrequest_from_sa :  STD_LOGIC;
                signal internal_pcp_cpu_data_master_granted_niosII_openMac_clock_3_in :  STD_LOGIC;
                signal internal_pcp_cpu_data_master_qualified_request_niosII_openMac_clock_3_in :  STD_LOGIC;
                signal internal_pcp_cpu_data_master_requests_niosII_openMac_clock_3_in :  STD_LOGIC;
                signal niosII_openMac_clock_3_in_allgrants :  STD_LOGIC;
                signal niosII_openMac_clock_3_in_allow_new_arb_cycle :  STD_LOGIC;
                signal niosII_openMac_clock_3_in_any_bursting_master_saved_grant :  STD_LOGIC;
                signal niosII_openMac_clock_3_in_any_continuerequest :  STD_LOGIC;
                signal niosII_openMac_clock_3_in_arb_counter_enable :  STD_LOGIC;
                signal niosII_openMac_clock_3_in_arb_share_counter :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal niosII_openMac_clock_3_in_arb_share_counter_next_value :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal niosII_openMac_clock_3_in_arb_share_set_values :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal niosII_openMac_clock_3_in_beginbursttransfer_internal :  STD_LOGIC;
                signal niosII_openMac_clock_3_in_begins_xfer :  STD_LOGIC;
                signal niosII_openMac_clock_3_in_end_xfer :  STD_LOGIC;
                signal niosII_openMac_clock_3_in_firsttransfer :  STD_LOGIC;
                signal niosII_openMac_clock_3_in_grant_vector :  STD_LOGIC;
                signal niosII_openMac_clock_3_in_in_a_read_cycle :  STD_LOGIC;
                signal niosII_openMac_clock_3_in_in_a_write_cycle :  STD_LOGIC;
                signal niosII_openMac_clock_3_in_master_qreq_vector :  STD_LOGIC;
                signal niosII_openMac_clock_3_in_non_bursting_master_requests :  STD_LOGIC;
                signal niosII_openMac_clock_3_in_reg_firsttransfer :  STD_LOGIC;
                signal niosII_openMac_clock_3_in_slavearbiterlockenable :  STD_LOGIC;
                signal niosII_openMac_clock_3_in_slavearbiterlockenable2 :  STD_LOGIC;
                signal niosII_openMac_clock_3_in_unreg_firsttransfer :  STD_LOGIC;
                signal niosII_openMac_clock_3_in_waits_for_read :  STD_LOGIC;
                signal niosII_openMac_clock_3_in_waits_for_write :  STD_LOGIC;
                signal pcp_cpu_data_master_arbiterlock :  STD_LOGIC;
                signal pcp_cpu_data_master_arbiterlock2 :  STD_LOGIC;
                signal pcp_cpu_data_master_continuerequest :  STD_LOGIC;
                signal pcp_cpu_data_master_saved_grant_niosII_openMac_clock_3_in :  STD_LOGIC;
                signal wait_for_niosII_openMac_clock_3_in_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT niosII_openMac_clock_3_in_end_xfer;
    end if;

  end process;

  niosII_openMac_clock_3_in_begins_xfer <= NOT d1_reasons_to_wait AND (internal_pcp_cpu_data_master_qualified_request_niosII_openMac_clock_3_in);
  --assign niosII_openMac_clock_3_in_readdata_from_sa = niosII_openMac_clock_3_in_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  niosII_openMac_clock_3_in_readdata_from_sa <= niosII_openMac_clock_3_in_readdata;
  internal_pcp_cpu_data_master_requests_niosII_openMac_clock_3_in <= to_std_logic(((Std_Logic_Vector'(pcp_cpu_data_master_address_to_slave(25 DOWNTO 4) & std_logic_vector'("0000")) = std_logic_vector'("00000000000000100100000000")))) AND ((pcp_cpu_data_master_read OR pcp_cpu_data_master_write));
  --assign niosII_openMac_clock_3_in_waitrequest_from_sa = niosII_openMac_clock_3_in_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_niosII_openMac_clock_3_in_waitrequest_from_sa <= niosII_openMac_clock_3_in_waitrequest;
  --niosII_openMac_clock_3_in_arb_share_counter set values, which is an e_mux
  niosII_openMac_clock_3_in_arb_share_set_values <= std_logic_vector'("01");
  --niosII_openMac_clock_3_in_non_bursting_master_requests mux, which is an e_mux
  niosII_openMac_clock_3_in_non_bursting_master_requests <= internal_pcp_cpu_data_master_requests_niosII_openMac_clock_3_in;
  --niosII_openMac_clock_3_in_any_bursting_master_saved_grant mux, which is an e_mux
  niosII_openMac_clock_3_in_any_bursting_master_saved_grant <= std_logic'('0');
  --niosII_openMac_clock_3_in_arb_share_counter_next_value assignment, which is an e_assign
  niosII_openMac_clock_3_in_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(niosII_openMac_clock_3_in_firsttransfer) = '1'), (((std_logic_vector'("0000000000000000000000000000000") & (niosII_openMac_clock_3_in_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(niosII_openMac_clock_3_in_arb_share_counter)) = '1'), (((std_logic_vector'("0000000000000000000000000000000") & (niosII_openMac_clock_3_in_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 2);
  --niosII_openMac_clock_3_in_allgrants all slave grants, which is an e_mux
  niosII_openMac_clock_3_in_allgrants <= niosII_openMac_clock_3_in_grant_vector;
  --niosII_openMac_clock_3_in_end_xfer assignment, which is an e_assign
  niosII_openMac_clock_3_in_end_xfer <= NOT ((niosII_openMac_clock_3_in_waits_for_read OR niosII_openMac_clock_3_in_waits_for_write));
  --end_xfer_arb_share_counter_term_niosII_openMac_clock_3_in arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_niosII_openMac_clock_3_in <= niosII_openMac_clock_3_in_end_xfer AND (((NOT niosII_openMac_clock_3_in_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --niosII_openMac_clock_3_in_arb_share_counter arbitration counter enable, which is an e_assign
  niosII_openMac_clock_3_in_arb_counter_enable <= ((end_xfer_arb_share_counter_term_niosII_openMac_clock_3_in AND niosII_openMac_clock_3_in_allgrants)) OR ((end_xfer_arb_share_counter_term_niosII_openMac_clock_3_in AND NOT niosII_openMac_clock_3_in_non_bursting_master_requests));
  --niosII_openMac_clock_3_in_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_openMac_clock_3_in_arb_share_counter <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      if std_logic'(niosII_openMac_clock_3_in_arb_counter_enable) = '1' then 
        niosII_openMac_clock_3_in_arb_share_counter <= niosII_openMac_clock_3_in_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --niosII_openMac_clock_3_in_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_openMac_clock_3_in_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((niosII_openMac_clock_3_in_master_qreq_vector AND end_xfer_arb_share_counter_term_niosII_openMac_clock_3_in)) OR ((end_xfer_arb_share_counter_term_niosII_openMac_clock_3_in AND NOT niosII_openMac_clock_3_in_non_bursting_master_requests)))) = '1' then 
        niosII_openMac_clock_3_in_slavearbiterlockenable <= or_reduce(niosII_openMac_clock_3_in_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --pcp_cpu/data_master niosII_openMac_clock_3/in arbiterlock, which is an e_assign
  pcp_cpu_data_master_arbiterlock <= niosII_openMac_clock_3_in_slavearbiterlockenable AND pcp_cpu_data_master_continuerequest;
  --niosII_openMac_clock_3_in_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  niosII_openMac_clock_3_in_slavearbiterlockenable2 <= or_reduce(niosII_openMac_clock_3_in_arb_share_counter_next_value);
  --pcp_cpu/data_master niosII_openMac_clock_3/in arbiterlock2, which is an e_assign
  pcp_cpu_data_master_arbiterlock2 <= niosII_openMac_clock_3_in_slavearbiterlockenable2 AND pcp_cpu_data_master_continuerequest;
  --niosII_openMac_clock_3_in_any_continuerequest at least one master continues requesting, which is an e_assign
  niosII_openMac_clock_3_in_any_continuerequest <= std_logic'('1');
  --pcp_cpu_data_master_continuerequest continued request, which is an e_assign
  pcp_cpu_data_master_continuerequest <= std_logic'('1');
  internal_pcp_cpu_data_master_qualified_request_niosII_openMac_clock_3_in <= internal_pcp_cpu_data_master_requests_niosII_openMac_clock_3_in AND NOT ((((pcp_cpu_data_master_read AND (NOT pcp_cpu_data_master_waitrequest))) OR (((NOT pcp_cpu_data_master_waitrequest) AND pcp_cpu_data_master_write))));
  --niosII_openMac_clock_3_in_writedata mux, which is an e_mux
  niosII_openMac_clock_3_in_writedata <= pcp_cpu_data_master_writedata;
  --assign niosII_openMac_clock_3_in_endofpacket_from_sa = niosII_openMac_clock_3_in_endofpacket so that symbol knows where to group signals which may go to master only, which is an e_assign
  niosII_openMac_clock_3_in_endofpacket_from_sa <= niosII_openMac_clock_3_in_endofpacket;
  --master is always granted when requested
  internal_pcp_cpu_data_master_granted_niosII_openMac_clock_3_in <= internal_pcp_cpu_data_master_qualified_request_niosII_openMac_clock_3_in;
  --pcp_cpu/data_master saved-grant niosII_openMac_clock_3/in, which is an e_assign
  pcp_cpu_data_master_saved_grant_niosII_openMac_clock_3_in <= internal_pcp_cpu_data_master_requests_niosII_openMac_clock_3_in;
  --allow new arb cycle for niosII_openMac_clock_3/in, which is an e_assign
  niosII_openMac_clock_3_in_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  niosII_openMac_clock_3_in_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  niosII_openMac_clock_3_in_master_qreq_vector <= std_logic'('1');
  --niosII_openMac_clock_3_in_reset_n assignment, which is an e_assign
  niosII_openMac_clock_3_in_reset_n <= reset_n;
  --niosII_openMac_clock_3_in_firsttransfer first transaction, which is an e_assign
  niosII_openMac_clock_3_in_firsttransfer <= A_WE_StdLogic((std_logic'(niosII_openMac_clock_3_in_begins_xfer) = '1'), niosII_openMac_clock_3_in_unreg_firsttransfer, niosII_openMac_clock_3_in_reg_firsttransfer);
  --niosII_openMac_clock_3_in_unreg_firsttransfer first transaction, which is an e_assign
  niosII_openMac_clock_3_in_unreg_firsttransfer <= NOT ((niosII_openMac_clock_3_in_slavearbiterlockenable AND niosII_openMac_clock_3_in_any_continuerequest));
  --niosII_openMac_clock_3_in_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_openMac_clock_3_in_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(niosII_openMac_clock_3_in_begins_xfer) = '1' then 
        niosII_openMac_clock_3_in_reg_firsttransfer <= niosII_openMac_clock_3_in_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --niosII_openMac_clock_3_in_beginbursttransfer_internal begin burst transfer, which is an e_assign
  niosII_openMac_clock_3_in_beginbursttransfer_internal <= niosII_openMac_clock_3_in_begins_xfer;
  --niosII_openMac_clock_3_in_read assignment, which is an e_mux
  niosII_openMac_clock_3_in_read <= internal_pcp_cpu_data_master_granted_niosII_openMac_clock_3_in AND pcp_cpu_data_master_read;
  --niosII_openMac_clock_3_in_write assignment, which is an e_mux
  niosII_openMac_clock_3_in_write <= internal_pcp_cpu_data_master_granted_niosII_openMac_clock_3_in AND pcp_cpu_data_master_write;
  --niosII_openMac_clock_3_in_address mux, which is an e_mux
  niosII_openMac_clock_3_in_address <= pcp_cpu_data_master_address_to_slave (3 DOWNTO 0);
  --slaveid niosII_openMac_clock_3_in_nativeaddress nativeaddress mux, which is an e_mux
  niosII_openMac_clock_3_in_nativeaddress <= A_EXT (A_SRL(pcp_cpu_data_master_address_to_slave,std_logic_vector'("00000000000000000000000000000010")), 2);
  --d1_niosII_openMac_clock_3_in_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_niosII_openMac_clock_3_in_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_niosII_openMac_clock_3_in_end_xfer <= niosII_openMac_clock_3_in_end_xfer;
    end if;

  end process;

  --niosII_openMac_clock_3_in_waits_for_read in a cycle, which is an e_mux
  niosII_openMac_clock_3_in_waits_for_read <= niosII_openMac_clock_3_in_in_a_read_cycle AND internal_niosII_openMac_clock_3_in_waitrequest_from_sa;
  --niosII_openMac_clock_3_in_in_a_read_cycle assignment, which is an e_assign
  niosII_openMac_clock_3_in_in_a_read_cycle <= internal_pcp_cpu_data_master_granted_niosII_openMac_clock_3_in AND pcp_cpu_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= niosII_openMac_clock_3_in_in_a_read_cycle;
  --niosII_openMac_clock_3_in_waits_for_write in a cycle, which is an e_mux
  niosII_openMac_clock_3_in_waits_for_write <= niosII_openMac_clock_3_in_in_a_write_cycle AND internal_niosII_openMac_clock_3_in_waitrequest_from_sa;
  --niosII_openMac_clock_3_in_in_a_write_cycle assignment, which is an e_assign
  niosII_openMac_clock_3_in_in_a_write_cycle <= internal_pcp_cpu_data_master_granted_niosII_openMac_clock_3_in AND pcp_cpu_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= niosII_openMac_clock_3_in_in_a_write_cycle;
  wait_for_niosII_openMac_clock_3_in_counter <= std_logic'('0');
  --niosII_openMac_clock_3_in_byteenable byte enable port mux, which is an e_mux
  niosII_openMac_clock_3_in_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_pcp_cpu_data_master_granted_niosII_openMac_clock_3_in)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (pcp_cpu_data_master_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))), 4);
  --vhdl renameroo for output signals
  niosII_openMac_clock_3_in_waitrequest_from_sa <= internal_niosII_openMac_clock_3_in_waitrequest_from_sa;
  --vhdl renameroo for output signals
  pcp_cpu_data_master_granted_niosII_openMac_clock_3_in <= internal_pcp_cpu_data_master_granted_niosII_openMac_clock_3_in;
  --vhdl renameroo for output signals
  pcp_cpu_data_master_qualified_request_niosII_openMac_clock_3_in <= internal_pcp_cpu_data_master_qualified_request_niosII_openMac_clock_3_in;
  --vhdl renameroo for output signals
  pcp_cpu_data_master_requests_niosII_openMac_clock_3_in <= internal_pcp_cpu_data_master_requests_niosII_openMac_clock_3_in;
--synthesis translate_off
    --niosII_openMac_clock_3/in enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity niosII_openMac_clock_3_out_arbitrator is 
        port (
              -- inputs:
                 signal altpll_0_pll_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal clk : IN STD_LOGIC;
                 signal d1_altpll_0_pll_slave_end_xfer : IN STD_LOGIC;
                 signal niosII_openMac_clock_3_out_address : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal niosII_openMac_clock_3_out_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal niosII_openMac_clock_3_out_granted_altpll_0_pll_slave : IN STD_LOGIC;
                 signal niosII_openMac_clock_3_out_qualified_request_altpll_0_pll_slave : IN STD_LOGIC;
                 signal niosII_openMac_clock_3_out_read : IN STD_LOGIC;
                 signal niosII_openMac_clock_3_out_read_data_valid_altpll_0_pll_slave : IN STD_LOGIC;
                 signal niosII_openMac_clock_3_out_requests_altpll_0_pll_slave : IN STD_LOGIC;
                 signal niosII_openMac_clock_3_out_write : IN STD_LOGIC;
                 signal niosII_openMac_clock_3_out_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal niosII_openMac_clock_3_out_address_to_slave : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal niosII_openMac_clock_3_out_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal niosII_openMac_clock_3_out_reset_n : OUT STD_LOGIC;
                 signal niosII_openMac_clock_3_out_waitrequest : OUT STD_LOGIC
              );
end entity niosII_openMac_clock_3_out_arbitrator;


architecture europa of niosII_openMac_clock_3_out_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal internal_niosII_openMac_clock_3_out_address_to_slave :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal internal_niosII_openMac_clock_3_out_waitrequest :  STD_LOGIC;
                signal niosII_openMac_clock_3_out_address_last_time :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_openMac_clock_3_out_byteenable_last_time :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_openMac_clock_3_out_read_last_time :  STD_LOGIC;
                signal niosII_openMac_clock_3_out_run :  STD_LOGIC;
                signal niosII_openMac_clock_3_out_write_last_time :  STD_LOGIC;
                signal niosII_openMac_clock_3_out_writedata_last_time :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal r_0 :  STD_LOGIC;

begin

  --r_0 master_run cascaded wait assignment, which is an e_assign
  r_0 <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000001") AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT niosII_openMac_clock_3_out_qualified_request_altpll_0_pll_slave OR NOT ((niosII_openMac_clock_3_out_read OR niosII_openMac_clock_3_out_write)))))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((niosII_openMac_clock_3_out_read OR niosII_openMac_clock_3_out_write)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT niosII_openMac_clock_3_out_qualified_request_altpll_0_pll_slave OR NOT ((niosII_openMac_clock_3_out_read OR niosII_openMac_clock_3_out_write)))))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((niosII_openMac_clock_3_out_read OR niosII_openMac_clock_3_out_write)))))))))));
  --cascaded wait assignment, which is an e_assign
  niosII_openMac_clock_3_out_run <= r_0;
  --optimize select-logic by passing only those address bits which matter.
  internal_niosII_openMac_clock_3_out_address_to_slave <= niosII_openMac_clock_3_out_address;
  --niosII_openMac_clock_3/out readdata mux, which is an e_mux
  niosII_openMac_clock_3_out_readdata <= altpll_0_pll_slave_readdata_from_sa;
  --actual waitrequest port, which is an e_assign
  internal_niosII_openMac_clock_3_out_waitrequest <= NOT niosII_openMac_clock_3_out_run;
  --niosII_openMac_clock_3_out_reset_n assignment, which is an e_assign
  niosII_openMac_clock_3_out_reset_n <= reset_n;
  --vhdl renameroo for output signals
  niosII_openMac_clock_3_out_address_to_slave <= internal_niosII_openMac_clock_3_out_address_to_slave;
  --vhdl renameroo for output signals
  niosII_openMac_clock_3_out_waitrequest <= internal_niosII_openMac_clock_3_out_waitrequest;
--synthesis translate_off
    --niosII_openMac_clock_3_out_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_openMac_clock_3_out_address_last_time <= std_logic_vector'("0000");
      elsif clk'event and clk = '1' then
        niosII_openMac_clock_3_out_address_last_time <= niosII_openMac_clock_3_out_address;
      end if;

    end process;

    --niosII_openMac_clock_3/out waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_niosII_openMac_clock_3_out_waitrequest AND ((niosII_openMac_clock_3_out_read OR niosII_openMac_clock_3_out_write));
      end if;

    end process;

    --niosII_openMac_clock_3_out_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line31 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((niosII_openMac_clock_3_out_address /= niosII_openMac_clock_3_out_address_last_time))))) = '1' then 
          write(write_line31, now);
          write(write_line31, string'(": "));
          write(write_line31, string'("niosII_openMac_clock_3_out_address did not heed wait!!!"));
          write(output, write_line31.all);
          deallocate (write_line31);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_openMac_clock_3_out_byteenable check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_openMac_clock_3_out_byteenable_last_time <= std_logic_vector'("0000");
      elsif clk'event and clk = '1' then
        niosII_openMac_clock_3_out_byteenable_last_time <= niosII_openMac_clock_3_out_byteenable;
      end if;

    end process;

    --niosII_openMac_clock_3_out_byteenable matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line32 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((niosII_openMac_clock_3_out_byteenable /= niosII_openMac_clock_3_out_byteenable_last_time))))) = '1' then 
          write(write_line32, now);
          write(write_line32, string'(": "));
          write(write_line32, string'("niosII_openMac_clock_3_out_byteenable did not heed wait!!!"));
          write(output, write_line32.all);
          deallocate (write_line32);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_openMac_clock_3_out_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_openMac_clock_3_out_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        niosII_openMac_clock_3_out_read_last_time <= niosII_openMac_clock_3_out_read;
      end if;

    end process;

    --niosII_openMac_clock_3_out_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line33 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(niosII_openMac_clock_3_out_read) /= std_logic'(niosII_openMac_clock_3_out_read_last_time)))))) = '1' then 
          write(write_line33, now);
          write(write_line33, string'(": "));
          write(write_line33, string'("niosII_openMac_clock_3_out_read did not heed wait!!!"));
          write(output, write_line33.all);
          deallocate (write_line33);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_openMac_clock_3_out_write check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_openMac_clock_3_out_write_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        niosII_openMac_clock_3_out_write_last_time <= niosII_openMac_clock_3_out_write;
      end if;

    end process;

    --niosII_openMac_clock_3_out_write matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line34 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(niosII_openMac_clock_3_out_write) /= std_logic'(niosII_openMac_clock_3_out_write_last_time)))))) = '1' then 
          write(write_line34, now);
          write(write_line34, string'(": "));
          write(write_line34, string'("niosII_openMac_clock_3_out_write did not heed wait!!!"));
          write(output, write_line34.all);
          deallocate (write_line34);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_openMac_clock_3_out_writedata check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_openMac_clock_3_out_writedata_last_time <= std_logic_vector'("00000000000000000000000000000000");
      elsif clk'event and clk = '1' then
        niosII_openMac_clock_3_out_writedata_last_time <= niosII_openMac_clock_3_out_writedata;
      end if;

    end process;

    --niosII_openMac_clock_3_out_writedata matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line35 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((active_and_waiting_last_time AND to_std_logic(((niosII_openMac_clock_3_out_writedata /= niosII_openMac_clock_3_out_writedata_last_time)))) AND niosII_openMac_clock_3_out_write)) = '1' then 
          write(write_line35, now);
          write(write_line35, string'(": "));
          write(write_line35, string'("niosII_openMac_clock_3_out_writedata did not heed wait!!!"));
          write(output, write_line35.all);
          deallocate (write_line35);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity niosII_openMac_clock_4_in_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal niosII_openMac_clock_4_in_endofpacket : IN STD_LOGIC;
                 signal niosII_openMac_clock_4_in_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal niosII_openMac_clock_4_in_waitrequest : IN STD_LOGIC;
                 signal pcp_cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (25 DOWNTO 0);
                 signal pcp_cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal pcp_cpu_data_master_read : IN STD_LOGIC;
                 signal pcp_cpu_data_master_waitrequest : IN STD_LOGIC;
                 signal pcp_cpu_data_master_write : IN STD_LOGIC;
                 signal pcp_cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal d1_niosII_openMac_clock_4_in_end_xfer : OUT STD_LOGIC;
                 signal niosII_openMac_clock_4_in_address : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal niosII_openMac_clock_4_in_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal niosII_openMac_clock_4_in_endofpacket_from_sa : OUT STD_LOGIC;
                 signal niosII_openMac_clock_4_in_nativeaddress : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
                 signal niosII_openMac_clock_4_in_read : OUT STD_LOGIC;
                 signal niosII_openMac_clock_4_in_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal niosII_openMac_clock_4_in_reset_n : OUT STD_LOGIC;
                 signal niosII_openMac_clock_4_in_waitrequest_from_sa : OUT STD_LOGIC;
                 signal niosII_openMac_clock_4_in_write : OUT STD_LOGIC;
                 signal niosII_openMac_clock_4_in_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal pcp_cpu_data_master_granted_niosII_openMac_clock_4_in : OUT STD_LOGIC;
                 signal pcp_cpu_data_master_qualified_request_niosII_openMac_clock_4_in : OUT STD_LOGIC;
                 signal pcp_cpu_data_master_read_data_valid_niosII_openMac_clock_4_in : OUT STD_LOGIC;
                 signal pcp_cpu_data_master_requests_niosII_openMac_clock_4_in : OUT STD_LOGIC
              );
end entity niosII_openMac_clock_4_in_arbitrator;


architecture europa of niosII_openMac_clock_4_in_arbitrator is
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_niosII_openMac_clock_4_in :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_niosII_openMac_clock_4_in_waitrequest_from_sa :  STD_LOGIC;
                signal internal_pcp_cpu_data_master_granted_niosII_openMac_clock_4_in :  STD_LOGIC;
                signal internal_pcp_cpu_data_master_qualified_request_niosII_openMac_clock_4_in :  STD_LOGIC;
                signal internal_pcp_cpu_data_master_requests_niosII_openMac_clock_4_in :  STD_LOGIC;
                signal niosII_openMac_clock_4_in_allgrants :  STD_LOGIC;
                signal niosII_openMac_clock_4_in_allow_new_arb_cycle :  STD_LOGIC;
                signal niosII_openMac_clock_4_in_any_bursting_master_saved_grant :  STD_LOGIC;
                signal niosII_openMac_clock_4_in_any_continuerequest :  STD_LOGIC;
                signal niosII_openMac_clock_4_in_arb_counter_enable :  STD_LOGIC;
                signal niosII_openMac_clock_4_in_arb_share_counter :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal niosII_openMac_clock_4_in_arb_share_counter_next_value :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal niosII_openMac_clock_4_in_arb_share_set_values :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal niosII_openMac_clock_4_in_beginbursttransfer_internal :  STD_LOGIC;
                signal niosII_openMac_clock_4_in_begins_xfer :  STD_LOGIC;
                signal niosII_openMac_clock_4_in_end_xfer :  STD_LOGIC;
                signal niosII_openMac_clock_4_in_firsttransfer :  STD_LOGIC;
                signal niosII_openMac_clock_4_in_grant_vector :  STD_LOGIC;
                signal niosII_openMac_clock_4_in_in_a_read_cycle :  STD_LOGIC;
                signal niosII_openMac_clock_4_in_in_a_write_cycle :  STD_LOGIC;
                signal niosII_openMac_clock_4_in_master_qreq_vector :  STD_LOGIC;
                signal niosII_openMac_clock_4_in_non_bursting_master_requests :  STD_LOGIC;
                signal niosII_openMac_clock_4_in_reg_firsttransfer :  STD_LOGIC;
                signal niosII_openMac_clock_4_in_slavearbiterlockenable :  STD_LOGIC;
                signal niosII_openMac_clock_4_in_slavearbiterlockenable2 :  STD_LOGIC;
                signal niosII_openMac_clock_4_in_unreg_firsttransfer :  STD_LOGIC;
                signal niosII_openMac_clock_4_in_waits_for_read :  STD_LOGIC;
                signal niosII_openMac_clock_4_in_waits_for_write :  STD_LOGIC;
                signal pcp_cpu_data_master_arbiterlock :  STD_LOGIC;
                signal pcp_cpu_data_master_arbiterlock2 :  STD_LOGIC;
                signal pcp_cpu_data_master_continuerequest :  STD_LOGIC;
                signal pcp_cpu_data_master_saved_grant_niosII_openMac_clock_4_in :  STD_LOGIC;
                signal shifted_address_to_niosII_openMac_clock_4_in_from_pcp_cpu_data_master :  STD_LOGIC_VECTOR (25 DOWNTO 0);
                signal wait_for_niosII_openMac_clock_4_in_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT niosII_openMac_clock_4_in_end_xfer;
    end if;

  end process;

  niosII_openMac_clock_4_in_begins_xfer <= NOT d1_reasons_to_wait AND (internal_pcp_cpu_data_master_qualified_request_niosII_openMac_clock_4_in);
  --assign niosII_openMac_clock_4_in_readdata_from_sa = niosII_openMac_clock_4_in_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  niosII_openMac_clock_4_in_readdata_from_sa <= niosII_openMac_clock_4_in_readdata;
  internal_pcp_cpu_data_master_requests_niosII_openMac_clock_4_in <= to_std_logic(((Std_Logic_Vector'(pcp_cpu_data_master_address_to_slave(25 DOWNTO 8) & std_logic_vector'("00000000")) = std_logic_vector'("00000000000000100000000000")))) AND ((pcp_cpu_data_master_read OR pcp_cpu_data_master_write));
  --assign niosII_openMac_clock_4_in_waitrequest_from_sa = niosII_openMac_clock_4_in_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_niosII_openMac_clock_4_in_waitrequest_from_sa <= niosII_openMac_clock_4_in_waitrequest;
  --niosII_openMac_clock_4_in_arb_share_counter set values, which is an e_mux
  niosII_openMac_clock_4_in_arb_share_set_values <= std_logic_vector'("01");
  --niosII_openMac_clock_4_in_non_bursting_master_requests mux, which is an e_mux
  niosII_openMac_clock_4_in_non_bursting_master_requests <= internal_pcp_cpu_data_master_requests_niosII_openMac_clock_4_in;
  --niosII_openMac_clock_4_in_any_bursting_master_saved_grant mux, which is an e_mux
  niosII_openMac_clock_4_in_any_bursting_master_saved_grant <= std_logic'('0');
  --niosII_openMac_clock_4_in_arb_share_counter_next_value assignment, which is an e_assign
  niosII_openMac_clock_4_in_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(niosII_openMac_clock_4_in_firsttransfer) = '1'), (((std_logic_vector'("0000000000000000000000000000000") & (niosII_openMac_clock_4_in_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(niosII_openMac_clock_4_in_arb_share_counter)) = '1'), (((std_logic_vector'("0000000000000000000000000000000") & (niosII_openMac_clock_4_in_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 2);
  --niosII_openMac_clock_4_in_allgrants all slave grants, which is an e_mux
  niosII_openMac_clock_4_in_allgrants <= niosII_openMac_clock_4_in_grant_vector;
  --niosII_openMac_clock_4_in_end_xfer assignment, which is an e_assign
  niosII_openMac_clock_4_in_end_xfer <= NOT ((niosII_openMac_clock_4_in_waits_for_read OR niosII_openMac_clock_4_in_waits_for_write));
  --end_xfer_arb_share_counter_term_niosII_openMac_clock_4_in arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_niosII_openMac_clock_4_in <= niosII_openMac_clock_4_in_end_xfer AND (((NOT niosII_openMac_clock_4_in_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --niosII_openMac_clock_4_in_arb_share_counter arbitration counter enable, which is an e_assign
  niosII_openMac_clock_4_in_arb_counter_enable <= ((end_xfer_arb_share_counter_term_niosII_openMac_clock_4_in AND niosII_openMac_clock_4_in_allgrants)) OR ((end_xfer_arb_share_counter_term_niosII_openMac_clock_4_in AND NOT niosII_openMac_clock_4_in_non_bursting_master_requests));
  --niosII_openMac_clock_4_in_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_openMac_clock_4_in_arb_share_counter <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      if std_logic'(niosII_openMac_clock_4_in_arb_counter_enable) = '1' then 
        niosII_openMac_clock_4_in_arb_share_counter <= niosII_openMac_clock_4_in_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --niosII_openMac_clock_4_in_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_openMac_clock_4_in_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((niosII_openMac_clock_4_in_master_qreq_vector AND end_xfer_arb_share_counter_term_niosII_openMac_clock_4_in)) OR ((end_xfer_arb_share_counter_term_niosII_openMac_clock_4_in AND NOT niosII_openMac_clock_4_in_non_bursting_master_requests)))) = '1' then 
        niosII_openMac_clock_4_in_slavearbiterlockenable <= or_reduce(niosII_openMac_clock_4_in_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --pcp_cpu/data_master niosII_openMac_clock_4/in arbiterlock, which is an e_assign
  pcp_cpu_data_master_arbiterlock <= niosII_openMac_clock_4_in_slavearbiterlockenable AND pcp_cpu_data_master_continuerequest;
  --niosII_openMac_clock_4_in_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  niosII_openMac_clock_4_in_slavearbiterlockenable2 <= or_reduce(niosII_openMac_clock_4_in_arb_share_counter_next_value);
  --pcp_cpu/data_master niosII_openMac_clock_4/in arbiterlock2, which is an e_assign
  pcp_cpu_data_master_arbiterlock2 <= niosII_openMac_clock_4_in_slavearbiterlockenable2 AND pcp_cpu_data_master_continuerequest;
  --niosII_openMac_clock_4_in_any_continuerequest at least one master continues requesting, which is an e_assign
  niosII_openMac_clock_4_in_any_continuerequest <= std_logic'('1');
  --pcp_cpu_data_master_continuerequest continued request, which is an e_assign
  pcp_cpu_data_master_continuerequest <= std_logic'('1');
  internal_pcp_cpu_data_master_qualified_request_niosII_openMac_clock_4_in <= internal_pcp_cpu_data_master_requests_niosII_openMac_clock_4_in AND NOT ((((pcp_cpu_data_master_read AND (NOT pcp_cpu_data_master_waitrequest))) OR (((NOT pcp_cpu_data_master_waitrequest) AND pcp_cpu_data_master_write))));
  --niosII_openMac_clock_4_in_writedata mux, which is an e_mux
  niosII_openMac_clock_4_in_writedata <= pcp_cpu_data_master_writedata;
  --assign niosII_openMac_clock_4_in_endofpacket_from_sa = niosII_openMac_clock_4_in_endofpacket so that symbol knows where to group signals which may go to master only, which is an e_assign
  niosII_openMac_clock_4_in_endofpacket_from_sa <= niosII_openMac_clock_4_in_endofpacket;
  --master is always granted when requested
  internal_pcp_cpu_data_master_granted_niosII_openMac_clock_4_in <= internal_pcp_cpu_data_master_qualified_request_niosII_openMac_clock_4_in;
  --pcp_cpu/data_master saved-grant niosII_openMac_clock_4/in, which is an e_assign
  pcp_cpu_data_master_saved_grant_niosII_openMac_clock_4_in <= internal_pcp_cpu_data_master_requests_niosII_openMac_clock_4_in;
  --allow new arb cycle for niosII_openMac_clock_4/in, which is an e_assign
  niosII_openMac_clock_4_in_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  niosII_openMac_clock_4_in_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  niosII_openMac_clock_4_in_master_qreq_vector <= std_logic'('1');
  --niosII_openMac_clock_4_in_reset_n assignment, which is an e_assign
  niosII_openMac_clock_4_in_reset_n <= reset_n;
  --niosII_openMac_clock_4_in_firsttransfer first transaction, which is an e_assign
  niosII_openMac_clock_4_in_firsttransfer <= A_WE_StdLogic((std_logic'(niosII_openMac_clock_4_in_begins_xfer) = '1'), niosII_openMac_clock_4_in_unreg_firsttransfer, niosII_openMac_clock_4_in_reg_firsttransfer);
  --niosII_openMac_clock_4_in_unreg_firsttransfer first transaction, which is an e_assign
  niosII_openMac_clock_4_in_unreg_firsttransfer <= NOT ((niosII_openMac_clock_4_in_slavearbiterlockenable AND niosII_openMac_clock_4_in_any_continuerequest));
  --niosII_openMac_clock_4_in_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_openMac_clock_4_in_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(niosII_openMac_clock_4_in_begins_xfer) = '1' then 
        niosII_openMac_clock_4_in_reg_firsttransfer <= niosII_openMac_clock_4_in_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --niosII_openMac_clock_4_in_beginbursttransfer_internal begin burst transfer, which is an e_assign
  niosII_openMac_clock_4_in_beginbursttransfer_internal <= niosII_openMac_clock_4_in_begins_xfer;
  --niosII_openMac_clock_4_in_read assignment, which is an e_mux
  niosII_openMac_clock_4_in_read <= internal_pcp_cpu_data_master_granted_niosII_openMac_clock_4_in AND pcp_cpu_data_master_read;
  --niosII_openMac_clock_4_in_write assignment, which is an e_mux
  niosII_openMac_clock_4_in_write <= internal_pcp_cpu_data_master_granted_niosII_openMac_clock_4_in AND pcp_cpu_data_master_write;
  shifted_address_to_niosII_openMac_clock_4_in_from_pcp_cpu_data_master <= pcp_cpu_data_master_address_to_slave;
  --niosII_openMac_clock_4_in_address mux, which is an e_mux
  niosII_openMac_clock_4_in_address <= A_EXT (A_SRL(shifted_address_to_niosII_openMac_clock_4_in_from_pcp_cpu_data_master,std_logic_vector'("00000000000000000000000000000010")), 8);
  --slaveid niosII_openMac_clock_4_in_nativeaddress nativeaddress mux, which is an e_mux
  niosII_openMac_clock_4_in_nativeaddress <= A_EXT (A_SRL(pcp_cpu_data_master_address_to_slave,std_logic_vector'("00000000000000000000000000000010")), 6);
  --d1_niosII_openMac_clock_4_in_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_niosII_openMac_clock_4_in_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_niosII_openMac_clock_4_in_end_xfer <= niosII_openMac_clock_4_in_end_xfer;
    end if;

  end process;

  --niosII_openMac_clock_4_in_waits_for_read in a cycle, which is an e_mux
  niosII_openMac_clock_4_in_waits_for_read <= niosII_openMac_clock_4_in_in_a_read_cycle AND internal_niosII_openMac_clock_4_in_waitrequest_from_sa;
  --niosII_openMac_clock_4_in_in_a_read_cycle assignment, which is an e_assign
  niosII_openMac_clock_4_in_in_a_read_cycle <= internal_pcp_cpu_data_master_granted_niosII_openMac_clock_4_in AND pcp_cpu_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= niosII_openMac_clock_4_in_in_a_read_cycle;
  --niosII_openMac_clock_4_in_waits_for_write in a cycle, which is an e_mux
  niosII_openMac_clock_4_in_waits_for_write <= niosII_openMac_clock_4_in_in_a_write_cycle AND internal_niosII_openMac_clock_4_in_waitrequest_from_sa;
  --niosII_openMac_clock_4_in_in_a_write_cycle assignment, which is an e_assign
  niosII_openMac_clock_4_in_in_a_write_cycle <= internal_pcp_cpu_data_master_granted_niosII_openMac_clock_4_in AND pcp_cpu_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= niosII_openMac_clock_4_in_in_a_write_cycle;
  wait_for_niosII_openMac_clock_4_in_counter <= std_logic'('0');
  --niosII_openMac_clock_4_in_byteenable byte enable port mux, which is an e_mux
  niosII_openMac_clock_4_in_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_pcp_cpu_data_master_granted_niosII_openMac_clock_4_in)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (pcp_cpu_data_master_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))), 4);
  --vhdl renameroo for output signals
  niosII_openMac_clock_4_in_waitrequest_from_sa <= internal_niosII_openMac_clock_4_in_waitrequest_from_sa;
  --vhdl renameroo for output signals
  pcp_cpu_data_master_granted_niosII_openMac_clock_4_in <= internal_pcp_cpu_data_master_granted_niosII_openMac_clock_4_in;
  --vhdl renameroo for output signals
  pcp_cpu_data_master_qualified_request_niosII_openMac_clock_4_in <= internal_pcp_cpu_data_master_qualified_request_niosII_openMac_clock_4_in;
  --vhdl renameroo for output signals
  pcp_cpu_data_master_requests_niosII_openMac_clock_4_in <= internal_pcp_cpu_data_master_requests_niosII_openMac_clock_4_in;
--synthesis translate_off
    --niosII_openMac_clock_4/in enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity niosII_openMac_clock_4_out_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal d1_remote_update_cycloneiii_0_s1_end_xfer : IN STD_LOGIC;
                 signal niosII_openMac_clock_4_out_address : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal niosII_openMac_clock_4_out_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal niosII_openMac_clock_4_out_granted_remote_update_cycloneiii_0_s1 : IN STD_LOGIC;
                 signal niosII_openMac_clock_4_out_qualified_request_remote_update_cycloneiii_0_s1 : IN STD_LOGIC;
                 signal niosII_openMac_clock_4_out_read : IN STD_LOGIC;
                 signal niosII_openMac_clock_4_out_read_data_valid_remote_update_cycloneiii_0_s1 : IN STD_LOGIC;
                 signal niosII_openMac_clock_4_out_requests_remote_update_cycloneiii_0_s1 : IN STD_LOGIC;
                 signal niosII_openMac_clock_4_out_write : IN STD_LOGIC;
                 signal niosII_openMac_clock_4_out_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal remote_update_cycloneiii_0_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal remote_update_cycloneiii_0_s1_waitrequest_from_sa : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal niosII_openMac_clock_4_out_address_to_slave : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal niosII_openMac_clock_4_out_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal niosII_openMac_clock_4_out_reset_n : OUT STD_LOGIC;
                 signal niosII_openMac_clock_4_out_waitrequest : OUT STD_LOGIC
              );
end entity niosII_openMac_clock_4_out_arbitrator;


architecture europa of niosII_openMac_clock_4_out_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal internal_niosII_openMac_clock_4_out_address_to_slave :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal internal_niosII_openMac_clock_4_out_waitrequest :  STD_LOGIC;
                signal niosII_openMac_clock_4_out_address_last_time :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal niosII_openMac_clock_4_out_byteenable_last_time :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_openMac_clock_4_out_read_last_time :  STD_LOGIC;
                signal niosII_openMac_clock_4_out_run :  STD_LOGIC;
                signal niosII_openMac_clock_4_out_write_last_time :  STD_LOGIC;
                signal niosII_openMac_clock_4_out_writedata_last_time :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal r_2 :  STD_LOGIC;

begin

  --r_2 master_run cascaded wait assignment, which is an e_assign
  r_2 <= Vector_To_Std_Logic((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((niosII_openMac_clock_4_out_qualified_request_remote_update_cycloneiii_0_s1 OR niosII_openMac_clock_4_out_read_data_valid_remote_update_cycloneiii_0_s1) OR NOT niosII_openMac_clock_4_out_requests_remote_update_cycloneiii_0_s1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((NOT niosII_openMac_clock_4_out_qualified_request_remote_update_cycloneiii_0_s1 OR NOT niosII_openMac_clock_4_out_read) OR ((niosII_openMac_clock_4_out_read_data_valid_remote_update_cycloneiii_0_s1 AND niosII_openMac_clock_4_out_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT niosII_openMac_clock_4_out_qualified_request_remote_update_cycloneiii_0_s1 OR NOT ((niosII_openMac_clock_4_out_read OR niosII_openMac_clock_4_out_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT remote_update_cycloneiii_0_s1_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((niosII_openMac_clock_4_out_read OR niosII_openMac_clock_4_out_write)))))))))));
  --cascaded wait assignment, which is an e_assign
  niosII_openMac_clock_4_out_run <= r_2;
  --optimize select-logic by passing only those address bits which matter.
  internal_niosII_openMac_clock_4_out_address_to_slave <= niosII_openMac_clock_4_out_address;
  --niosII_openMac_clock_4/out readdata mux, which is an e_mux
  niosII_openMac_clock_4_out_readdata <= remote_update_cycloneiii_0_s1_readdata_from_sa;
  --actual waitrequest port, which is an e_assign
  internal_niosII_openMac_clock_4_out_waitrequest <= NOT niosII_openMac_clock_4_out_run;
  --niosII_openMac_clock_4_out_reset_n assignment, which is an e_assign
  niosII_openMac_clock_4_out_reset_n <= reset_n;
  --vhdl renameroo for output signals
  niosII_openMac_clock_4_out_address_to_slave <= internal_niosII_openMac_clock_4_out_address_to_slave;
  --vhdl renameroo for output signals
  niosII_openMac_clock_4_out_waitrequest <= internal_niosII_openMac_clock_4_out_waitrequest;
--synthesis translate_off
    --niosII_openMac_clock_4_out_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_openMac_clock_4_out_address_last_time <= std_logic_vector'("00000000");
      elsif clk'event and clk = '1' then
        niosII_openMac_clock_4_out_address_last_time <= niosII_openMac_clock_4_out_address;
      end if;

    end process;

    --niosII_openMac_clock_4/out waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_niosII_openMac_clock_4_out_waitrequest AND ((niosII_openMac_clock_4_out_read OR niosII_openMac_clock_4_out_write));
      end if;

    end process;

    --niosII_openMac_clock_4_out_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line36 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((niosII_openMac_clock_4_out_address /= niosII_openMac_clock_4_out_address_last_time))))) = '1' then 
          write(write_line36, now);
          write(write_line36, string'(": "));
          write(write_line36, string'("niosII_openMac_clock_4_out_address did not heed wait!!!"));
          write(output, write_line36.all);
          deallocate (write_line36);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_openMac_clock_4_out_byteenable check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_openMac_clock_4_out_byteenable_last_time <= std_logic_vector'("0000");
      elsif clk'event and clk = '1' then
        niosII_openMac_clock_4_out_byteenable_last_time <= niosII_openMac_clock_4_out_byteenable;
      end if;

    end process;

    --niosII_openMac_clock_4_out_byteenable matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line37 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((niosII_openMac_clock_4_out_byteenable /= niosII_openMac_clock_4_out_byteenable_last_time))))) = '1' then 
          write(write_line37, now);
          write(write_line37, string'(": "));
          write(write_line37, string'("niosII_openMac_clock_4_out_byteenable did not heed wait!!!"));
          write(output, write_line37.all);
          deallocate (write_line37);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_openMac_clock_4_out_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_openMac_clock_4_out_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        niosII_openMac_clock_4_out_read_last_time <= niosII_openMac_clock_4_out_read;
      end if;

    end process;

    --niosII_openMac_clock_4_out_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line38 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(niosII_openMac_clock_4_out_read) /= std_logic'(niosII_openMac_clock_4_out_read_last_time)))))) = '1' then 
          write(write_line38, now);
          write(write_line38, string'(": "));
          write(write_line38, string'("niosII_openMac_clock_4_out_read did not heed wait!!!"));
          write(output, write_line38.all);
          deallocate (write_line38);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_openMac_clock_4_out_write check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_openMac_clock_4_out_write_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        niosII_openMac_clock_4_out_write_last_time <= niosII_openMac_clock_4_out_write;
      end if;

    end process;

    --niosII_openMac_clock_4_out_write matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line39 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(niosII_openMac_clock_4_out_write) /= std_logic'(niosII_openMac_clock_4_out_write_last_time)))))) = '1' then 
          write(write_line39, now);
          write(write_line39, string'(": "));
          write(write_line39, string'("niosII_openMac_clock_4_out_write did not heed wait!!!"));
          write(output, write_line39.all);
          deallocate (write_line39);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --niosII_openMac_clock_4_out_writedata check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        niosII_openMac_clock_4_out_writedata_last_time <= std_logic_vector'("00000000000000000000000000000000");
      elsif clk'event and clk = '1' then
        niosII_openMac_clock_4_out_writedata_last_time <= niosII_openMac_clock_4_out_writedata;
      end if;

    end process;

    --niosII_openMac_clock_4_out_writedata matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line40 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((active_and_waiting_last_time AND to_std_logic(((niosII_openMac_clock_4_out_writedata /= niosII_openMac_clock_4_out_writedata_last_time)))) AND niosII_openMac_clock_4_out_write)) = '1' then 
          write(write_line40, now);
          write(write_line40, string'(": "));
          write(write_line40, string'("niosII_openMac_clock_4_out_writedata did not heed wait!!!"));
          write(output, write_line40.all);
          deallocate (write_line40);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity node_switch_pio_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal clock_crossing_1_m1_address_to_slave : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal clock_crossing_1_m1_latency_counter : IN STD_LOGIC;
                 signal clock_crossing_1_m1_nativeaddress : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
                 signal clock_crossing_1_m1_read : IN STD_LOGIC;
                 signal clock_crossing_1_m1_write : IN STD_LOGIC;
                 signal node_switch_pio_s1_readdata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal clock_crossing_1_m1_granted_node_switch_pio_s1 : OUT STD_LOGIC;
                 signal clock_crossing_1_m1_qualified_request_node_switch_pio_s1 : OUT STD_LOGIC;
                 signal clock_crossing_1_m1_read_data_valid_node_switch_pio_s1 : OUT STD_LOGIC;
                 signal clock_crossing_1_m1_requests_node_switch_pio_s1 : OUT STD_LOGIC;
                 signal d1_node_switch_pio_s1_end_xfer : OUT STD_LOGIC;
                 signal node_switch_pio_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal node_switch_pio_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal node_switch_pio_s1_reset_n : OUT STD_LOGIC
              );
end entity node_switch_pio_s1_arbitrator;


architecture europa of node_switch_pio_s1_arbitrator is
                signal clock_crossing_1_m1_arbiterlock :  STD_LOGIC;
                signal clock_crossing_1_m1_arbiterlock2 :  STD_LOGIC;
                signal clock_crossing_1_m1_continuerequest :  STD_LOGIC;
                signal clock_crossing_1_m1_saved_grant_node_switch_pio_s1 :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_node_switch_pio_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_clock_crossing_1_m1_granted_node_switch_pio_s1 :  STD_LOGIC;
                signal internal_clock_crossing_1_m1_qualified_request_node_switch_pio_s1 :  STD_LOGIC;
                signal internal_clock_crossing_1_m1_requests_node_switch_pio_s1 :  STD_LOGIC;
                signal node_switch_pio_s1_allgrants :  STD_LOGIC;
                signal node_switch_pio_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal node_switch_pio_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal node_switch_pio_s1_any_continuerequest :  STD_LOGIC;
                signal node_switch_pio_s1_arb_counter_enable :  STD_LOGIC;
                signal node_switch_pio_s1_arb_share_counter :  STD_LOGIC;
                signal node_switch_pio_s1_arb_share_counter_next_value :  STD_LOGIC;
                signal node_switch_pio_s1_arb_share_set_values :  STD_LOGIC;
                signal node_switch_pio_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal node_switch_pio_s1_begins_xfer :  STD_LOGIC;
                signal node_switch_pio_s1_end_xfer :  STD_LOGIC;
                signal node_switch_pio_s1_firsttransfer :  STD_LOGIC;
                signal node_switch_pio_s1_grant_vector :  STD_LOGIC;
                signal node_switch_pio_s1_in_a_read_cycle :  STD_LOGIC;
                signal node_switch_pio_s1_in_a_write_cycle :  STD_LOGIC;
                signal node_switch_pio_s1_master_qreq_vector :  STD_LOGIC;
                signal node_switch_pio_s1_non_bursting_master_requests :  STD_LOGIC;
                signal node_switch_pio_s1_reg_firsttransfer :  STD_LOGIC;
                signal node_switch_pio_s1_slavearbiterlockenable :  STD_LOGIC;
                signal node_switch_pio_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal node_switch_pio_s1_unreg_firsttransfer :  STD_LOGIC;
                signal node_switch_pio_s1_waits_for_read :  STD_LOGIC;
                signal node_switch_pio_s1_waits_for_write :  STD_LOGIC;
                signal wait_for_node_switch_pio_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT node_switch_pio_s1_end_xfer;
    end if;

  end process;

  node_switch_pio_s1_begins_xfer <= NOT d1_reasons_to_wait AND (internal_clock_crossing_1_m1_qualified_request_node_switch_pio_s1);
  --assign node_switch_pio_s1_readdata_from_sa = node_switch_pio_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  node_switch_pio_s1_readdata_from_sa <= node_switch_pio_s1_readdata;
  internal_clock_crossing_1_m1_requests_node_switch_pio_s1 <= ((to_std_logic(((Std_Logic_Vector'(clock_crossing_1_m1_address_to_slave(7 DOWNTO 4) & std_logic_vector'("0000")) = std_logic_vector'("10110000")))) AND ((clock_crossing_1_m1_read OR clock_crossing_1_m1_write)))) AND clock_crossing_1_m1_read;
  --node_switch_pio_s1_arb_share_counter set values, which is an e_mux
  node_switch_pio_s1_arb_share_set_values <= std_logic'('1');
  --node_switch_pio_s1_non_bursting_master_requests mux, which is an e_mux
  node_switch_pio_s1_non_bursting_master_requests <= internal_clock_crossing_1_m1_requests_node_switch_pio_s1;
  --node_switch_pio_s1_any_bursting_master_saved_grant mux, which is an e_mux
  node_switch_pio_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --node_switch_pio_s1_arb_share_counter_next_value assignment, which is an e_assign
  node_switch_pio_s1_arb_share_counter_next_value <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(node_switch_pio_s1_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(node_switch_pio_s1_arb_share_set_values))) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(node_switch_pio_s1_arb_share_counter) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(node_switch_pio_s1_arb_share_counter))) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))));
  --node_switch_pio_s1_allgrants all slave grants, which is an e_mux
  node_switch_pio_s1_allgrants <= node_switch_pio_s1_grant_vector;
  --node_switch_pio_s1_end_xfer assignment, which is an e_assign
  node_switch_pio_s1_end_xfer <= NOT ((node_switch_pio_s1_waits_for_read OR node_switch_pio_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_node_switch_pio_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_node_switch_pio_s1 <= node_switch_pio_s1_end_xfer AND (((NOT node_switch_pio_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --node_switch_pio_s1_arb_share_counter arbitration counter enable, which is an e_assign
  node_switch_pio_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_node_switch_pio_s1 AND node_switch_pio_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_node_switch_pio_s1 AND NOT node_switch_pio_s1_non_bursting_master_requests));
  --node_switch_pio_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      node_switch_pio_s1_arb_share_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(node_switch_pio_s1_arb_counter_enable) = '1' then 
        node_switch_pio_s1_arb_share_counter <= node_switch_pio_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --node_switch_pio_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      node_switch_pio_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((node_switch_pio_s1_master_qreq_vector AND end_xfer_arb_share_counter_term_node_switch_pio_s1)) OR ((end_xfer_arb_share_counter_term_node_switch_pio_s1 AND NOT node_switch_pio_s1_non_bursting_master_requests)))) = '1' then 
        node_switch_pio_s1_slavearbiterlockenable <= node_switch_pio_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --clock_crossing_1/m1 node_switch_pio/s1 arbiterlock, which is an e_assign
  clock_crossing_1_m1_arbiterlock <= node_switch_pio_s1_slavearbiterlockenable AND clock_crossing_1_m1_continuerequest;
  --node_switch_pio_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  node_switch_pio_s1_slavearbiterlockenable2 <= node_switch_pio_s1_arb_share_counter_next_value;
  --clock_crossing_1/m1 node_switch_pio/s1 arbiterlock2, which is an e_assign
  clock_crossing_1_m1_arbiterlock2 <= node_switch_pio_s1_slavearbiterlockenable2 AND clock_crossing_1_m1_continuerequest;
  --node_switch_pio_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  node_switch_pio_s1_any_continuerequest <= std_logic'('1');
  --clock_crossing_1_m1_continuerequest continued request, which is an e_assign
  clock_crossing_1_m1_continuerequest <= std_logic'('1');
  internal_clock_crossing_1_m1_qualified_request_node_switch_pio_s1 <= internal_clock_crossing_1_m1_requests_node_switch_pio_s1 AND NOT ((clock_crossing_1_m1_read AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(clock_crossing_1_m1_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))))));
  --local readdatavalid clock_crossing_1_m1_read_data_valid_node_switch_pio_s1, which is an e_mux
  clock_crossing_1_m1_read_data_valid_node_switch_pio_s1 <= (internal_clock_crossing_1_m1_granted_node_switch_pio_s1 AND clock_crossing_1_m1_read) AND NOT node_switch_pio_s1_waits_for_read;
  --master is always granted when requested
  internal_clock_crossing_1_m1_granted_node_switch_pio_s1 <= internal_clock_crossing_1_m1_qualified_request_node_switch_pio_s1;
  --clock_crossing_1/m1 saved-grant node_switch_pio/s1, which is an e_assign
  clock_crossing_1_m1_saved_grant_node_switch_pio_s1 <= internal_clock_crossing_1_m1_requests_node_switch_pio_s1;
  --allow new arb cycle for node_switch_pio/s1, which is an e_assign
  node_switch_pio_s1_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  node_switch_pio_s1_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  node_switch_pio_s1_master_qreq_vector <= std_logic'('1');
  --node_switch_pio_s1_reset_n assignment, which is an e_assign
  node_switch_pio_s1_reset_n <= reset_n;
  --node_switch_pio_s1_firsttransfer first transaction, which is an e_assign
  node_switch_pio_s1_firsttransfer <= A_WE_StdLogic((std_logic'(node_switch_pio_s1_begins_xfer) = '1'), node_switch_pio_s1_unreg_firsttransfer, node_switch_pio_s1_reg_firsttransfer);
  --node_switch_pio_s1_unreg_firsttransfer first transaction, which is an e_assign
  node_switch_pio_s1_unreg_firsttransfer <= NOT ((node_switch_pio_s1_slavearbiterlockenable AND node_switch_pio_s1_any_continuerequest));
  --node_switch_pio_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      node_switch_pio_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(node_switch_pio_s1_begins_xfer) = '1' then 
        node_switch_pio_s1_reg_firsttransfer <= node_switch_pio_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --node_switch_pio_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  node_switch_pio_s1_beginbursttransfer_internal <= node_switch_pio_s1_begins_xfer;
  --node_switch_pio_s1_address mux, which is an e_mux
  node_switch_pio_s1_address <= clock_crossing_1_m1_nativeaddress (1 DOWNTO 0);
  --d1_node_switch_pio_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_node_switch_pio_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_node_switch_pio_s1_end_xfer <= node_switch_pio_s1_end_xfer;
    end if;

  end process;

  --node_switch_pio_s1_waits_for_read in a cycle, which is an e_mux
  node_switch_pio_s1_waits_for_read <= node_switch_pio_s1_in_a_read_cycle AND node_switch_pio_s1_begins_xfer;
  --node_switch_pio_s1_in_a_read_cycle assignment, which is an e_assign
  node_switch_pio_s1_in_a_read_cycle <= internal_clock_crossing_1_m1_granted_node_switch_pio_s1 AND clock_crossing_1_m1_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= node_switch_pio_s1_in_a_read_cycle;
  --node_switch_pio_s1_waits_for_write in a cycle, which is an e_mux
  node_switch_pio_s1_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(node_switch_pio_s1_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --node_switch_pio_s1_in_a_write_cycle assignment, which is an e_assign
  node_switch_pio_s1_in_a_write_cycle <= internal_clock_crossing_1_m1_granted_node_switch_pio_s1 AND clock_crossing_1_m1_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= node_switch_pio_s1_in_a_write_cycle;
  wait_for_node_switch_pio_s1_counter <= std_logic'('0');
  --vhdl renameroo for output signals
  clock_crossing_1_m1_granted_node_switch_pio_s1 <= internal_clock_crossing_1_m1_granted_node_switch_pio_s1;
  --vhdl renameroo for output signals
  clock_crossing_1_m1_qualified_request_node_switch_pio_s1 <= internal_clock_crossing_1_m1_qualified_request_node_switch_pio_s1;
  --vhdl renameroo for output signals
  clock_crossing_1_m1_requests_node_switch_pio_s1 <= internal_clock_crossing_1_m1_requests_node_switch_pio_s1;
--synthesis translate_off
    --node_switch_pio/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity onchip_memory_0_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal onchip_memory_0_s1_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal pcp_cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (25 DOWNTO 0);
                 signal pcp_cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal pcp_cpu_data_master_read : IN STD_LOGIC;
                 signal pcp_cpu_data_master_waitrequest : IN STD_LOGIC;
                 signal pcp_cpu_data_master_write : IN STD_LOGIC;
                 signal pcp_cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal pcp_cpu_instruction_master_address_to_slave : IN STD_LOGIC_VECTOR (25 DOWNTO 0);
                 signal pcp_cpu_instruction_master_latency_counter : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal pcp_cpu_instruction_master_read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal d1_onchip_memory_0_s1_end_xfer : OUT STD_LOGIC;
                 signal onchip_memory_0_s1_address : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal onchip_memory_0_s1_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal onchip_memory_0_s1_chipselect : OUT STD_LOGIC;
                 signal onchip_memory_0_s1_clken : OUT STD_LOGIC;
                 signal onchip_memory_0_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal onchip_memory_0_s1_write : OUT STD_LOGIC;
                 signal onchip_memory_0_s1_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal pcp_cpu_data_master_granted_onchip_memory_0_s1 : OUT STD_LOGIC;
                 signal pcp_cpu_data_master_qualified_request_onchip_memory_0_s1 : OUT STD_LOGIC;
                 signal pcp_cpu_data_master_read_data_valid_onchip_memory_0_s1 : OUT STD_LOGIC;
                 signal pcp_cpu_data_master_requests_onchip_memory_0_s1 : OUT STD_LOGIC;
                 signal pcp_cpu_instruction_master_granted_onchip_memory_0_s1 : OUT STD_LOGIC;
                 signal pcp_cpu_instruction_master_qualified_request_onchip_memory_0_s1 : OUT STD_LOGIC;
                 signal pcp_cpu_instruction_master_read_data_valid_onchip_memory_0_s1 : OUT STD_LOGIC;
                 signal pcp_cpu_instruction_master_requests_onchip_memory_0_s1 : OUT STD_LOGIC;
                 signal registered_pcp_cpu_data_master_read_data_valid_onchip_memory_0_s1 : OUT STD_LOGIC
              );
end entity onchip_memory_0_s1_arbitrator;


architecture europa of onchip_memory_0_s1_arbitrator is
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_onchip_memory_0_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_pcp_cpu_data_master_granted_onchip_memory_0_s1 :  STD_LOGIC;
                signal internal_pcp_cpu_data_master_qualified_request_onchip_memory_0_s1 :  STD_LOGIC;
                signal internal_pcp_cpu_data_master_requests_onchip_memory_0_s1 :  STD_LOGIC;
                signal internal_pcp_cpu_instruction_master_granted_onchip_memory_0_s1 :  STD_LOGIC;
                signal internal_pcp_cpu_instruction_master_qualified_request_onchip_memory_0_s1 :  STD_LOGIC;
                signal internal_pcp_cpu_instruction_master_requests_onchip_memory_0_s1 :  STD_LOGIC;
                signal last_cycle_pcp_cpu_data_master_granted_slave_onchip_memory_0_s1 :  STD_LOGIC;
                signal last_cycle_pcp_cpu_instruction_master_granted_slave_onchip_memory_0_s1 :  STD_LOGIC;
                signal onchip_memory_0_s1_allgrants :  STD_LOGIC;
                signal onchip_memory_0_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal onchip_memory_0_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal onchip_memory_0_s1_any_continuerequest :  STD_LOGIC;
                signal onchip_memory_0_s1_arb_addend :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal onchip_memory_0_s1_arb_counter_enable :  STD_LOGIC;
                signal onchip_memory_0_s1_arb_share_counter :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal onchip_memory_0_s1_arb_share_counter_next_value :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal onchip_memory_0_s1_arb_share_set_values :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal onchip_memory_0_s1_arb_winner :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal onchip_memory_0_s1_arbitration_holdoff_internal :  STD_LOGIC;
                signal onchip_memory_0_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal onchip_memory_0_s1_begins_xfer :  STD_LOGIC;
                signal onchip_memory_0_s1_chosen_master_double_vector :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal onchip_memory_0_s1_chosen_master_rot_left :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal onchip_memory_0_s1_end_xfer :  STD_LOGIC;
                signal onchip_memory_0_s1_firsttransfer :  STD_LOGIC;
                signal onchip_memory_0_s1_grant_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal onchip_memory_0_s1_in_a_read_cycle :  STD_LOGIC;
                signal onchip_memory_0_s1_in_a_write_cycle :  STD_LOGIC;
                signal onchip_memory_0_s1_master_qreq_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal onchip_memory_0_s1_non_bursting_master_requests :  STD_LOGIC;
                signal onchip_memory_0_s1_reg_firsttransfer :  STD_LOGIC;
                signal onchip_memory_0_s1_saved_chosen_master_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal onchip_memory_0_s1_slavearbiterlockenable :  STD_LOGIC;
                signal onchip_memory_0_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal onchip_memory_0_s1_unreg_firsttransfer :  STD_LOGIC;
                signal onchip_memory_0_s1_waits_for_read :  STD_LOGIC;
                signal onchip_memory_0_s1_waits_for_write :  STD_LOGIC;
                signal p1_pcp_cpu_data_master_read_data_valid_onchip_memory_0_s1_shift_register :  STD_LOGIC;
                signal p1_pcp_cpu_instruction_master_read_data_valid_onchip_memory_0_s1_shift_register :  STD_LOGIC;
                signal pcp_cpu_data_master_arbiterlock :  STD_LOGIC;
                signal pcp_cpu_data_master_arbiterlock2 :  STD_LOGIC;
                signal pcp_cpu_data_master_continuerequest :  STD_LOGIC;
                signal pcp_cpu_data_master_read_data_valid_onchip_memory_0_s1_shift_register :  STD_LOGIC;
                signal pcp_cpu_data_master_read_data_valid_onchip_memory_0_s1_shift_register_in :  STD_LOGIC;
                signal pcp_cpu_data_master_saved_grant_onchip_memory_0_s1 :  STD_LOGIC;
                signal pcp_cpu_instruction_master_arbiterlock :  STD_LOGIC;
                signal pcp_cpu_instruction_master_arbiterlock2 :  STD_LOGIC;
                signal pcp_cpu_instruction_master_continuerequest :  STD_LOGIC;
                signal pcp_cpu_instruction_master_read_data_valid_onchip_memory_0_s1_shift_register :  STD_LOGIC;
                signal pcp_cpu_instruction_master_read_data_valid_onchip_memory_0_s1_shift_register_in :  STD_LOGIC;
                signal pcp_cpu_instruction_master_saved_grant_onchip_memory_0_s1 :  STD_LOGIC;
                signal shifted_address_to_onchip_memory_0_s1_from_pcp_cpu_data_master :  STD_LOGIC_VECTOR (25 DOWNTO 0);
                signal shifted_address_to_onchip_memory_0_s1_from_pcp_cpu_instruction_master :  STD_LOGIC_VECTOR (25 DOWNTO 0);
                signal wait_for_onchip_memory_0_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT onchip_memory_0_s1_end_xfer;
    end if;

  end process;

  onchip_memory_0_s1_begins_xfer <= NOT d1_reasons_to_wait AND ((internal_pcp_cpu_data_master_qualified_request_onchip_memory_0_s1 OR internal_pcp_cpu_instruction_master_qualified_request_onchip_memory_0_s1));
  --assign onchip_memory_0_s1_readdata_from_sa = onchip_memory_0_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  onchip_memory_0_s1_readdata_from_sa <= onchip_memory_0_s1_readdata;
  internal_pcp_cpu_data_master_requests_onchip_memory_0_s1 <= to_std_logic(((Std_Logic_Vector'(pcp_cpu_data_master_address_to_slave(25 DOWNTO 10) & std_logic_vector'("0000000000")) = std_logic_vector'("00000000000100000000000000")))) AND ((pcp_cpu_data_master_read OR pcp_cpu_data_master_write));
  --registered rdv signal_name registered_pcp_cpu_data_master_read_data_valid_onchip_memory_0_s1 assignment, which is an e_assign
  registered_pcp_cpu_data_master_read_data_valid_onchip_memory_0_s1 <= pcp_cpu_data_master_read_data_valid_onchip_memory_0_s1_shift_register_in;
  --onchip_memory_0_s1_arb_share_counter set values, which is an e_mux
  onchip_memory_0_s1_arb_share_set_values <= std_logic_vector'("01");
  --onchip_memory_0_s1_non_bursting_master_requests mux, which is an e_mux
  onchip_memory_0_s1_non_bursting_master_requests <= ((internal_pcp_cpu_data_master_requests_onchip_memory_0_s1 OR internal_pcp_cpu_instruction_master_requests_onchip_memory_0_s1) OR internal_pcp_cpu_data_master_requests_onchip_memory_0_s1) OR internal_pcp_cpu_instruction_master_requests_onchip_memory_0_s1;
  --onchip_memory_0_s1_any_bursting_master_saved_grant mux, which is an e_mux
  onchip_memory_0_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --onchip_memory_0_s1_arb_share_counter_next_value assignment, which is an e_assign
  onchip_memory_0_s1_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(onchip_memory_0_s1_firsttransfer) = '1'), (((std_logic_vector'("0000000000000000000000000000000") & (onchip_memory_0_s1_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(onchip_memory_0_s1_arb_share_counter)) = '1'), (((std_logic_vector'("0000000000000000000000000000000") & (onchip_memory_0_s1_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 2);
  --onchip_memory_0_s1_allgrants all slave grants, which is an e_mux
  onchip_memory_0_s1_allgrants <= (((or_reduce(onchip_memory_0_s1_grant_vector)) OR (or_reduce(onchip_memory_0_s1_grant_vector))) OR (or_reduce(onchip_memory_0_s1_grant_vector))) OR (or_reduce(onchip_memory_0_s1_grant_vector));
  --onchip_memory_0_s1_end_xfer assignment, which is an e_assign
  onchip_memory_0_s1_end_xfer <= NOT ((onchip_memory_0_s1_waits_for_read OR onchip_memory_0_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_onchip_memory_0_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_onchip_memory_0_s1 <= onchip_memory_0_s1_end_xfer AND (((NOT onchip_memory_0_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --onchip_memory_0_s1_arb_share_counter arbitration counter enable, which is an e_assign
  onchip_memory_0_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_onchip_memory_0_s1 AND onchip_memory_0_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_onchip_memory_0_s1 AND NOT onchip_memory_0_s1_non_bursting_master_requests));
  --onchip_memory_0_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      onchip_memory_0_s1_arb_share_counter <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      if std_logic'(onchip_memory_0_s1_arb_counter_enable) = '1' then 
        onchip_memory_0_s1_arb_share_counter <= onchip_memory_0_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --onchip_memory_0_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      onchip_memory_0_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((or_reduce(onchip_memory_0_s1_master_qreq_vector) AND end_xfer_arb_share_counter_term_onchip_memory_0_s1)) OR ((end_xfer_arb_share_counter_term_onchip_memory_0_s1 AND NOT onchip_memory_0_s1_non_bursting_master_requests)))) = '1' then 
        onchip_memory_0_s1_slavearbiterlockenable <= or_reduce(onchip_memory_0_s1_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --pcp_cpu/data_master onchip_memory_0/s1 arbiterlock, which is an e_assign
  pcp_cpu_data_master_arbiterlock <= onchip_memory_0_s1_slavearbiterlockenable AND pcp_cpu_data_master_continuerequest;
  --onchip_memory_0_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  onchip_memory_0_s1_slavearbiterlockenable2 <= or_reduce(onchip_memory_0_s1_arb_share_counter_next_value);
  --pcp_cpu/data_master onchip_memory_0/s1 arbiterlock2, which is an e_assign
  pcp_cpu_data_master_arbiterlock2 <= onchip_memory_0_s1_slavearbiterlockenable2 AND pcp_cpu_data_master_continuerequest;
  --pcp_cpu/instruction_master onchip_memory_0/s1 arbiterlock, which is an e_assign
  pcp_cpu_instruction_master_arbiterlock <= onchip_memory_0_s1_slavearbiterlockenable AND pcp_cpu_instruction_master_continuerequest;
  --pcp_cpu/instruction_master onchip_memory_0/s1 arbiterlock2, which is an e_assign
  pcp_cpu_instruction_master_arbiterlock2 <= onchip_memory_0_s1_slavearbiterlockenable2 AND pcp_cpu_instruction_master_continuerequest;
  --pcp_cpu/instruction_master granted onchip_memory_0/s1 last time, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      last_cycle_pcp_cpu_instruction_master_granted_slave_onchip_memory_0_s1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      last_cycle_pcp_cpu_instruction_master_granted_slave_onchip_memory_0_s1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(pcp_cpu_instruction_master_saved_grant_onchip_memory_0_s1) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((onchip_memory_0_s1_arbitration_holdoff_internal OR NOT internal_pcp_cpu_instruction_master_requests_onchip_memory_0_s1))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_pcp_cpu_instruction_master_granted_slave_onchip_memory_0_s1))))));
    end if;

  end process;

  --pcp_cpu_instruction_master_continuerequest continued request, which is an e_mux
  pcp_cpu_instruction_master_continuerequest <= last_cycle_pcp_cpu_instruction_master_granted_slave_onchip_memory_0_s1 AND internal_pcp_cpu_instruction_master_requests_onchip_memory_0_s1;
  --onchip_memory_0_s1_any_continuerequest at least one master continues requesting, which is an e_mux
  onchip_memory_0_s1_any_continuerequest <= pcp_cpu_instruction_master_continuerequest OR pcp_cpu_data_master_continuerequest;
  internal_pcp_cpu_data_master_qualified_request_onchip_memory_0_s1 <= internal_pcp_cpu_data_master_requests_onchip_memory_0_s1 AND NOT (((((pcp_cpu_data_master_read AND (pcp_cpu_data_master_read_data_valid_onchip_memory_0_s1_shift_register))) OR (((NOT pcp_cpu_data_master_waitrequest) AND pcp_cpu_data_master_write))) OR pcp_cpu_instruction_master_arbiterlock));
  --pcp_cpu_data_master_read_data_valid_onchip_memory_0_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  pcp_cpu_data_master_read_data_valid_onchip_memory_0_s1_shift_register_in <= ((internal_pcp_cpu_data_master_granted_onchip_memory_0_s1 AND pcp_cpu_data_master_read) AND NOT onchip_memory_0_s1_waits_for_read) AND NOT (pcp_cpu_data_master_read_data_valid_onchip_memory_0_s1_shift_register);
  --shift register p1 pcp_cpu_data_master_read_data_valid_onchip_memory_0_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  p1_pcp_cpu_data_master_read_data_valid_onchip_memory_0_s1_shift_register <= Vector_To_Std_Logic(Std_Logic_Vector'(A_ToStdLogicVector(pcp_cpu_data_master_read_data_valid_onchip_memory_0_s1_shift_register) & A_ToStdLogicVector(pcp_cpu_data_master_read_data_valid_onchip_memory_0_s1_shift_register_in)));
  --pcp_cpu_data_master_read_data_valid_onchip_memory_0_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pcp_cpu_data_master_read_data_valid_onchip_memory_0_s1_shift_register <= std_logic'('0');
    elsif clk'event and clk = '1' then
      pcp_cpu_data_master_read_data_valid_onchip_memory_0_s1_shift_register <= p1_pcp_cpu_data_master_read_data_valid_onchip_memory_0_s1_shift_register;
    end if;

  end process;

  --local readdatavalid pcp_cpu_data_master_read_data_valid_onchip_memory_0_s1, which is an e_mux
  pcp_cpu_data_master_read_data_valid_onchip_memory_0_s1 <= pcp_cpu_data_master_read_data_valid_onchip_memory_0_s1_shift_register;
  --onchip_memory_0_s1_writedata mux, which is an e_mux
  onchip_memory_0_s1_writedata <= pcp_cpu_data_master_writedata;
  --mux onchip_memory_0_s1_clken, which is an e_mux
  onchip_memory_0_s1_clken <= std_logic'('1');
  internal_pcp_cpu_instruction_master_requests_onchip_memory_0_s1 <= ((to_std_logic(((Std_Logic_Vector'(pcp_cpu_instruction_master_address_to_slave(25 DOWNTO 10) & std_logic_vector'("0000000000")) = std_logic_vector'("00000000000100000000000000")))) AND (pcp_cpu_instruction_master_read))) AND pcp_cpu_instruction_master_read;
  --pcp_cpu/data_master granted onchip_memory_0/s1 last time, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      last_cycle_pcp_cpu_data_master_granted_slave_onchip_memory_0_s1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      last_cycle_pcp_cpu_data_master_granted_slave_onchip_memory_0_s1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(pcp_cpu_data_master_saved_grant_onchip_memory_0_s1) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((onchip_memory_0_s1_arbitration_holdoff_internal OR NOT internal_pcp_cpu_data_master_requests_onchip_memory_0_s1))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_pcp_cpu_data_master_granted_slave_onchip_memory_0_s1))))));
    end if;

  end process;

  --pcp_cpu_data_master_continuerequest continued request, which is an e_mux
  pcp_cpu_data_master_continuerequest <= last_cycle_pcp_cpu_data_master_granted_slave_onchip_memory_0_s1 AND internal_pcp_cpu_data_master_requests_onchip_memory_0_s1;
  internal_pcp_cpu_instruction_master_qualified_request_onchip_memory_0_s1 <= internal_pcp_cpu_instruction_master_requests_onchip_memory_0_s1 AND NOT ((((pcp_cpu_instruction_master_read AND to_std_logic(((std_logic_vector'("00000000000000000000000000000001")<(std_logic_vector'("000000000000000000000000000000") & (pcp_cpu_instruction_master_latency_counter))))))) OR pcp_cpu_data_master_arbiterlock));
  --pcp_cpu_instruction_master_read_data_valid_onchip_memory_0_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  pcp_cpu_instruction_master_read_data_valid_onchip_memory_0_s1_shift_register_in <= (internal_pcp_cpu_instruction_master_granted_onchip_memory_0_s1 AND pcp_cpu_instruction_master_read) AND NOT onchip_memory_0_s1_waits_for_read;
  --shift register p1 pcp_cpu_instruction_master_read_data_valid_onchip_memory_0_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  p1_pcp_cpu_instruction_master_read_data_valid_onchip_memory_0_s1_shift_register <= Vector_To_Std_Logic(Std_Logic_Vector'(A_ToStdLogicVector(pcp_cpu_instruction_master_read_data_valid_onchip_memory_0_s1_shift_register) & A_ToStdLogicVector(pcp_cpu_instruction_master_read_data_valid_onchip_memory_0_s1_shift_register_in)));
  --pcp_cpu_instruction_master_read_data_valid_onchip_memory_0_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pcp_cpu_instruction_master_read_data_valid_onchip_memory_0_s1_shift_register <= std_logic'('0');
    elsif clk'event and clk = '1' then
      pcp_cpu_instruction_master_read_data_valid_onchip_memory_0_s1_shift_register <= p1_pcp_cpu_instruction_master_read_data_valid_onchip_memory_0_s1_shift_register;
    end if;

  end process;

  --local readdatavalid pcp_cpu_instruction_master_read_data_valid_onchip_memory_0_s1, which is an e_mux
  pcp_cpu_instruction_master_read_data_valid_onchip_memory_0_s1 <= pcp_cpu_instruction_master_read_data_valid_onchip_memory_0_s1_shift_register;
  --allow new arb cycle for onchip_memory_0/s1, which is an e_assign
  onchip_memory_0_s1_allow_new_arb_cycle <= NOT pcp_cpu_data_master_arbiterlock AND NOT pcp_cpu_instruction_master_arbiterlock;
  --pcp_cpu/instruction_master assignment into master qualified-requests vector for onchip_memory_0/s1, which is an e_assign
  onchip_memory_0_s1_master_qreq_vector(0) <= internal_pcp_cpu_instruction_master_qualified_request_onchip_memory_0_s1;
  --pcp_cpu/instruction_master grant onchip_memory_0/s1, which is an e_assign
  internal_pcp_cpu_instruction_master_granted_onchip_memory_0_s1 <= onchip_memory_0_s1_grant_vector(0);
  --pcp_cpu/instruction_master saved-grant onchip_memory_0/s1, which is an e_assign
  pcp_cpu_instruction_master_saved_grant_onchip_memory_0_s1 <= onchip_memory_0_s1_arb_winner(0) AND internal_pcp_cpu_instruction_master_requests_onchip_memory_0_s1;
  --pcp_cpu/data_master assignment into master qualified-requests vector for onchip_memory_0/s1, which is an e_assign
  onchip_memory_0_s1_master_qreq_vector(1) <= internal_pcp_cpu_data_master_qualified_request_onchip_memory_0_s1;
  --pcp_cpu/data_master grant onchip_memory_0/s1, which is an e_assign
  internal_pcp_cpu_data_master_granted_onchip_memory_0_s1 <= onchip_memory_0_s1_grant_vector(1);
  --pcp_cpu/data_master saved-grant onchip_memory_0/s1, which is an e_assign
  pcp_cpu_data_master_saved_grant_onchip_memory_0_s1 <= onchip_memory_0_s1_arb_winner(1) AND internal_pcp_cpu_data_master_requests_onchip_memory_0_s1;
  --onchip_memory_0/s1 chosen-master double-vector, which is an e_assign
  onchip_memory_0_s1_chosen_master_double_vector <= A_EXT (((std_logic_vector'("0") & ((onchip_memory_0_s1_master_qreq_vector & onchip_memory_0_s1_master_qreq_vector))) AND (((std_logic_vector'("0") & (Std_Logic_Vector'(NOT onchip_memory_0_s1_master_qreq_vector & NOT onchip_memory_0_s1_master_qreq_vector))) + (std_logic_vector'("000") & (onchip_memory_0_s1_arb_addend))))), 4);
  --stable onehot encoding of arb winner
  onchip_memory_0_s1_arb_winner <= A_WE_StdLogicVector((std_logic'(((onchip_memory_0_s1_allow_new_arb_cycle AND or_reduce(onchip_memory_0_s1_grant_vector)))) = '1'), onchip_memory_0_s1_grant_vector, onchip_memory_0_s1_saved_chosen_master_vector);
  --saved onchip_memory_0_s1_grant_vector, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      onchip_memory_0_s1_saved_chosen_master_vector <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      if std_logic'(onchip_memory_0_s1_allow_new_arb_cycle) = '1' then 
        onchip_memory_0_s1_saved_chosen_master_vector <= A_WE_StdLogicVector((std_logic'(or_reduce(onchip_memory_0_s1_grant_vector)) = '1'), onchip_memory_0_s1_grant_vector, onchip_memory_0_s1_saved_chosen_master_vector);
      end if;
    end if;

  end process;

  --onehot encoding of chosen master
  onchip_memory_0_s1_grant_vector <= Std_Logic_Vector'(A_ToStdLogicVector(((onchip_memory_0_s1_chosen_master_double_vector(1) OR onchip_memory_0_s1_chosen_master_double_vector(3)))) & A_ToStdLogicVector(((onchip_memory_0_s1_chosen_master_double_vector(0) OR onchip_memory_0_s1_chosen_master_double_vector(2)))));
  --onchip_memory_0/s1 chosen master rotated left, which is an e_assign
  onchip_memory_0_s1_chosen_master_rot_left <= A_EXT (A_WE_StdLogicVector((((A_SLL(onchip_memory_0_s1_arb_winner,std_logic_vector'("00000000000000000000000000000001")))) /= std_logic_vector'("00")), (std_logic_vector'("000000000000000000000000000000") & ((A_SLL(onchip_memory_0_s1_arb_winner,std_logic_vector'("00000000000000000000000000000001"))))), std_logic_vector'("00000000000000000000000000000001")), 2);
  --onchip_memory_0/s1's addend for next-master-grant
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      onchip_memory_0_s1_arb_addend <= std_logic_vector'("01");
    elsif clk'event and clk = '1' then
      if std_logic'(or_reduce(onchip_memory_0_s1_grant_vector)) = '1' then 
        onchip_memory_0_s1_arb_addend <= A_WE_StdLogicVector((std_logic'(onchip_memory_0_s1_end_xfer) = '1'), onchip_memory_0_s1_chosen_master_rot_left, onchip_memory_0_s1_grant_vector);
      end if;
    end if;

  end process;

  onchip_memory_0_s1_chipselect <= internal_pcp_cpu_data_master_granted_onchip_memory_0_s1 OR internal_pcp_cpu_instruction_master_granted_onchip_memory_0_s1;
  --onchip_memory_0_s1_firsttransfer first transaction, which is an e_assign
  onchip_memory_0_s1_firsttransfer <= A_WE_StdLogic((std_logic'(onchip_memory_0_s1_begins_xfer) = '1'), onchip_memory_0_s1_unreg_firsttransfer, onchip_memory_0_s1_reg_firsttransfer);
  --onchip_memory_0_s1_unreg_firsttransfer first transaction, which is an e_assign
  onchip_memory_0_s1_unreg_firsttransfer <= NOT ((onchip_memory_0_s1_slavearbiterlockenable AND onchip_memory_0_s1_any_continuerequest));
  --onchip_memory_0_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      onchip_memory_0_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(onchip_memory_0_s1_begins_xfer) = '1' then 
        onchip_memory_0_s1_reg_firsttransfer <= onchip_memory_0_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --onchip_memory_0_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  onchip_memory_0_s1_beginbursttransfer_internal <= onchip_memory_0_s1_begins_xfer;
  --onchip_memory_0_s1_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  onchip_memory_0_s1_arbitration_holdoff_internal <= onchip_memory_0_s1_begins_xfer AND onchip_memory_0_s1_firsttransfer;
  --onchip_memory_0_s1_write assignment, which is an e_mux
  onchip_memory_0_s1_write <= internal_pcp_cpu_data_master_granted_onchip_memory_0_s1 AND pcp_cpu_data_master_write;
  shifted_address_to_onchip_memory_0_s1_from_pcp_cpu_data_master <= pcp_cpu_data_master_address_to_slave;
  --onchip_memory_0_s1_address mux, which is an e_mux
  onchip_memory_0_s1_address <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_pcp_cpu_data_master_granted_onchip_memory_0_s1)) = '1'), (A_SRL(shifted_address_to_onchip_memory_0_s1_from_pcp_cpu_data_master,std_logic_vector'("00000000000000000000000000000010"))), (A_SRL(shifted_address_to_onchip_memory_0_s1_from_pcp_cpu_instruction_master,std_logic_vector'("00000000000000000000000000000010")))), 8);
  shifted_address_to_onchip_memory_0_s1_from_pcp_cpu_instruction_master <= pcp_cpu_instruction_master_address_to_slave;
  --d1_onchip_memory_0_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_onchip_memory_0_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_onchip_memory_0_s1_end_xfer <= onchip_memory_0_s1_end_xfer;
    end if;

  end process;

  --onchip_memory_0_s1_waits_for_read in a cycle, which is an e_mux
  onchip_memory_0_s1_waits_for_read <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(onchip_memory_0_s1_in_a_read_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --onchip_memory_0_s1_in_a_read_cycle assignment, which is an e_assign
  onchip_memory_0_s1_in_a_read_cycle <= ((internal_pcp_cpu_data_master_granted_onchip_memory_0_s1 AND pcp_cpu_data_master_read)) OR ((internal_pcp_cpu_instruction_master_granted_onchip_memory_0_s1 AND pcp_cpu_instruction_master_read));
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= onchip_memory_0_s1_in_a_read_cycle;
  --onchip_memory_0_s1_waits_for_write in a cycle, which is an e_mux
  onchip_memory_0_s1_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(onchip_memory_0_s1_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --onchip_memory_0_s1_in_a_write_cycle assignment, which is an e_assign
  onchip_memory_0_s1_in_a_write_cycle <= internal_pcp_cpu_data_master_granted_onchip_memory_0_s1 AND pcp_cpu_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= onchip_memory_0_s1_in_a_write_cycle;
  wait_for_onchip_memory_0_s1_counter <= std_logic'('0');
  --onchip_memory_0_s1_byteenable byte enable port mux, which is an e_mux
  onchip_memory_0_s1_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_pcp_cpu_data_master_granted_onchip_memory_0_s1)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (pcp_cpu_data_master_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))), 4);
  --vhdl renameroo for output signals
  pcp_cpu_data_master_granted_onchip_memory_0_s1 <= internal_pcp_cpu_data_master_granted_onchip_memory_0_s1;
  --vhdl renameroo for output signals
  pcp_cpu_data_master_qualified_request_onchip_memory_0_s1 <= internal_pcp_cpu_data_master_qualified_request_onchip_memory_0_s1;
  --vhdl renameroo for output signals
  pcp_cpu_data_master_requests_onchip_memory_0_s1 <= internal_pcp_cpu_data_master_requests_onchip_memory_0_s1;
  --vhdl renameroo for output signals
  pcp_cpu_instruction_master_granted_onchip_memory_0_s1 <= internal_pcp_cpu_instruction_master_granted_onchip_memory_0_s1;
  --vhdl renameroo for output signals
  pcp_cpu_instruction_master_qualified_request_onchip_memory_0_s1 <= internal_pcp_cpu_instruction_master_qualified_request_onchip_memory_0_s1;
  --vhdl renameroo for output signals
  pcp_cpu_instruction_master_requests_onchip_memory_0_s1 <= internal_pcp_cpu_instruction_master_requests_onchip_memory_0_s1;
--synthesis translate_off
    --onchip_memory_0/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --grant signals are active simultaneously, which is an e_process
    process (clk)
    VARIABLE write_line41 : line;
    begin
      if clk'event and clk = '1' then
        if (std_logic_vector'("000000000000000000000000000000") & (((std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(internal_pcp_cpu_data_master_granted_onchip_memory_0_s1))) + (std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(internal_pcp_cpu_instruction_master_granted_onchip_memory_0_s1))))))>std_logic_vector'("00000000000000000000000000000001") then 
          write(write_line41, now);
          write(write_line41, string'(": "));
          write(write_line41, string'("> 1 of grant signals are active simultaneously"));
          write(output, write_line41.all);
          deallocate (write_line41);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --saved_grant signals are active simultaneously, which is an e_process
    process (clk)
    VARIABLE write_line42 : line;
    begin
      if clk'event and clk = '1' then
        if (std_logic_vector'("000000000000000000000000000000") & (((std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(pcp_cpu_data_master_saved_grant_onchip_memory_0_s1))) + (std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(pcp_cpu_instruction_master_saved_grant_onchip_memory_0_s1))))))>std_logic_vector'("00000000000000000000000000000001") then 
          write(write_line42, now);
          write(write_line42, string'(": "));
          write(write_line42, string'("> 1 of saved_grant signals are active simultaneously"));
          write(output, write_line42.all);
          deallocate (write_line42);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity pcp_cpu_jtag_debug_module_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal pcp_cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (25 DOWNTO 0);
                 signal pcp_cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal pcp_cpu_data_master_debugaccess : IN STD_LOGIC;
                 signal pcp_cpu_data_master_read : IN STD_LOGIC;
                 signal pcp_cpu_data_master_waitrequest : IN STD_LOGIC;
                 signal pcp_cpu_data_master_write : IN STD_LOGIC;
                 signal pcp_cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal pcp_cpu_instruction_master_address_to_slave : IN STD_LOGIC_VECTOR (25 DOWNTO 0);
                 signal pcp_cpu_instruction_master_latency_counter : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal pcp_cpu_instruction_master_read : IN STD_LOGIC;
                 signal pcp_cpu_jtag_debug_module_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal pcp_cpu_jtag_debug_module_resetrequest : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal d1_pcp_cpu_jtag_debug_module_end_xfer : OUT STD_LOGIC;
                 signal pcp_cpu_data_master_granted_pcp_cpu_jtag_debug_module : OUT STD_LOGIC;
                 signal pcp_cpu_data_master_qualified_request_pcp_cpu_jtag_debug_module : OUT STD_LOGIC;
                 signal pcp_cpu_data_master_read_data_valid_pcp_cpu_jtag_debug_module : OUT STD_LOGIC;
                 signal pcp_cpu_data_master_requests_pcp_cpu_jtag_debug_module : OUT STD_LOGIC;
                 signal pcp_cpu_instruction_master_granted_pcp_cpu_jtag_debug_module : OUT STD_LOGIC;
                 signal pcp_cpu_instruction_master_qualified_request_pcp_cpu_jtag_debug_module : OUT STD_LOGIC;
                 signal pcp_cpu_instruction_master_read_data_valid_pcp_cpu_jtag_debug_module : OUT STD_LOGIC;
                 signal pcp_cpu_instruction_master_requests_pcp_cpu_jtag_debug_module : OUT STD_LOGIC;
                 signal pcp_cpu_jtag_debug_module_address : OUT STD_LOGIC_VECTOR (8 DOWNTO 0);
                 signal pcp_cpu_jtag_debug_module_begintransfer : OUT STD_LOGIC;
                 signal pcp_cpu_jtag_debug_module_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal pcp_cpu_jtag_debug_module_chipselect : OUT STD_LOGIC;
                 signal pcp_cpu_jtag_debug_module_debugaccess : OUT STD_LOGIC;
                 signal pcp_cpu_jtag_debug_module_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal pcp_cpu_jtag_debug_module_reset_n : OUT STD_LOGIC;
                 signal pcp_cpu_jtag_debug_module_resetrequest_from_sa : OUT STD_LOGIC;
                 signal pcp_cpu_jtag_debug_module_write : OUT STD_LOGIC;
                 signal pcp_cpu_jtag_debug_module_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
              );
end entity pcp_cpu_jtag_debug_module_arbitrator;


architecture europa of pcp_cpu_jtag_debug_module_arbitrator is
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_pcp_cpu_jtag_debug_module :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_pcp_cpu_data_master_granted_pcp_cpu_jtag_debug_module :  STD_LOGIC;
                signal internal_pcp_cpu_data_master_qualified_request_pcp_cpu_jtag_debug_module :  STD_LOGIC;
                signal internal_pcp_cpu_data_master_requests_pcp_cpu_jtag_debug_module :  STD_LOGIC;
                signal internal_pcp_cpu_instruction_master_granted_pcp_cpu_jtag_debug_module :  STD_LOGIC;
                signal internal_pcp_cpu_instruction_master_qualified_request_pcp_cpu_jtag_debug_module :  STD_LOGIC;
                signal internal_pcp_cpu_instruction_master_requests_pcp_cpu_jtag_debug_module :  STD_LOGIC;
                signal last_cycle_pcp_cpu_data_master_granted_slave_pcp_cpu_jtag_debug_module :  STD_LOGIC;
                signal last_cycle_pcp_cpu_instruction_master_granted_slave_pcp_cpu_jtag_debug_module :  STD_LOGIC;
                signal pcp_cpu_data_master_arbiterlock :  STD_LOGIC;
                signal pcp_cpu_data_master_arbiterlock2 :  STD_LOGIC;
                signal pcp_cpu_data_master_continuerequest :  STD_LOGIC;
                signal pcp_cpu_data_master_saved_grant_pcp_cpu_jtag_debug_module :  STD_LOGIC;
                signal pcp_cpu_instruction_master_arbiterlock :  STD_LOGIC;
                signal pcp_cpu_instruction_master_arbiterlock2 :  STD_LOGIC;
                signal pcp_cpu_instruction_master_continuerequest :  STD_LOGIC;
                signal pcp_cpu_instruction_master_saved_grant_pcp_cpu_jtag_debug_module :  STD_LOGIC;
                signal pcp_cpu_jtag_debug_module_allgrants :  STD_LOGIC;
                signal pcp_cpu_jtag_debug_module_allow_new_arb_cycle :  STD_LOGIC;
                signal pcp_cpu_jtag_debug_module_any_bursting_master_saved_grant :  STD_LOGIC;
                signal pcp_cpu_jtag_debug_module_any_continuerequest :  STD_LOGIC;
                signal pcp_cpu_jtag_debug_module_arb_addend :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal pcp_cpu_jtag_debug_module_arb_counter_enable :  STD_LOGIC;
                signal pcp_cpu_jtag_debug_module_arb_share_counter :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal pcp_cpu_jtag_debug_module_arb_share_counter_next_value :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal pcp_cpu_jtag_debug_module_arb_share_set_values :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal pcp_cpu_jtag_debug_module_arb_winner :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal pcp_cpu_jtag_debug_module_arbitration_holdoff_internal :  STD_LOGIC;
                signal pcp_cpu_jtag_debug_module_beginbursttransfer_internal :  STD_LOGIC;
                signal pcp_cpu_jtag_debug_module_begins_xfer :  STD_LOGIC;
                signal pcp_cpu_jtag_debug_module_chosen_master_double_vector :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal pcp_cpu_jtag_debug_module_chosen_master_rot_left :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal pcp_cpu_jtag_debug_module_end_xfer :  STD_LOGIC;
                signal pcp_cpu_jtag_debug_module_firsttransfer :  STD_LOGIC;
                signal pcp_cpu_jtag_debug_module_grant_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal pcp_cpu_jtag_debug_module_in_a_read_cycle :  STD_LOGIC;
                signal pcp_cpu_jtag_debug_module_in_a_write_cycle :  STD_LOGIC;
                signal pcp_cpu_jtag_debug_module_master_qreq_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal pcp_cpu_jtag_debug_module_non_bursting_master_requests :  STD_LOGIC;
                signal pcp_cpu_jtag_debug_module_reg_firsttransfer :  STD_LOGIC;
                signal pcp_cpu_jtag_debug_module_saved_chosen_master_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal pcp_cpu_jtag_debug_module_slavearbiterlockenable :  STD_LOGIC;
                signal pcp_cpu_jtag_debug_module_slavearbiterlockenable2 :  STD_LOGIC;
                signal pcp_cpu_jtag_debug_module_unreg_firsttransfer :  STD_LOGIC;
                signal pcp_cpu_jtag_debug_module_waits_for_read :  STD_LOGIC;
                signal pcp_cpu_jtag_debug_module_waits_for_write :  STD_LOGIC;
                signal shifted_address_to_pcp_cpu_jtag_debug_module_from_pcp_cpu_data_master :  STD_LOGIC_VECTOR (25 DOWNTO 0);
                signal shifted_address_to_pcp_cpu_jtag_debug_module_from_pcp_cpu_instruction_master :  STD_LOGIC_VECTOR (25 DOWNTO 0);
                signal wait_for_pcp_cpu_jtag_debug_module_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT pcp_cpu_jtag_debug_module_end_xfer;
    end if;

  end process;

  pcp_cpu_jtag_debug_module_begins_xfer <= NOT d1_reasons_to_wait AND ((internal_pcp_cpu_data_master_qualified_request_pcp_cpu_jtag_debug_module OR internal_pcp_cpu_instruction_master_qualified_request_pcp_cpu_jtag_debug_module));
  --assign pcp_cpu_jtag_debug_module_readdata_from_sa = pcp_cpu_jtag_debug_module_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  pcp_cpu_jtag_debug_module_readdata_from_sa <= pcp_cpu_jtag_debug_module_readdata;
  internal_pcp_cpu_data_master_requests_pcp_cpu_jtag_debug_module <= to_std_logic(((Std_Logic_Vector'(pcp_cpu_data_master_address_to_slave(25 DOWNTO 11) & std_logic_vector'("00000000000")) = std_logic_vector'("00000000000001100000000000")))) AND ((pcp_cpu_data_master_read OR pcp_cpu_data_master_write));
  --pcp_cpu_jtag_debug_module_arb_share_counter set values, which is an e_mux
  pcp_cpu_jtag_debug_module_arb_share_set_values <= std_logic_vector'("01");
  --pcp_cpu_jtag_debug_module_non_bursting_master_requests mux, which is an e_mux
  pcp_cpu_jtag_debug_module_non_bursting_master_requests <= ((internal_pcp_cpu_data_master_requests_pcp_cpu_jtag_debug_module OR internal_pcp_cpu_instruction_master_requests_pcp_cpu_jtag_debug_module) OR internal_pcp_cpu_data_master_requests_pcp_cpu_jtag_debug_module) OR internal_pcp_cpu_instruction_master_requests_pcp_cpu_jtag_debug_module;
  --pcp_cpu_jtag_debug_module_any_bursting_master_saved_grant mux, which is an e_mux
  pcp_cpu_jtag_debug_module_any_bursting_master_saved_grant <= std_logic'('0');
  --pcp_cpu_jtag_debug_module_arb_share_counter_next_value assignment, which is an e_assign
  pcp_cpu_jtag_debug_module_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(pcp_cpu_jtag_debug_module_firsttransfer) = '1'), (((std_logic_vector'("0000000000000000000000000000000") & (pcp_cpu_jtag_debug_module_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(pcp_cpu_jtag_debug_module_arb_share_counter)) = '1'), (((std_logic_vector'("0000000000000000000000000000000") & (pcp_cpu_jtag_debug_module_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 2);
  --pcp_cpu_jtag_debug_module_allgrants all slave grants, which is an e_mux
  pcp_cpu_jtag_debug_module_allgrants <= (((or_reduce(pcp_cpu_jtag_debug_module_grant_vector)) OR (or_reduce(pcp_cpu_jtag_debug_module_grant_vector))) OR (or_reduce(pcp_cpu_jtag_debug_module_grant_vector))) OR (or_reduce(pcp_cpu_jtag_debug_module_grant_vector));
  --pcp_cpu_jtag_debug_module_end_xfer assignment, which is an e_assign
  pcp_cpu_jtag_debug_module_end_xfer <= NOT ((pcp_cpu_jtag_debug_module_waits_for_read OR pcp_cpu_jtag_debug_module_waits_for_write));
  --end_xfer_arb_share_counter_term_pcp_cpu_jtag_debug_module arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_pcp_cpu_jtag_debug_module <= pcp_cpu_jtag_debug_module_end_xfer AND (((NOT pcp_cpu_jtag_debug_module_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --pcp_cpu_jtag_debug_module_arb_share_counter arbitration counter enable, which is an e_assign
  pcp_cpu_jtag_debug_module_arb_counter_enable <= ((end_xfer_arb_share_counter_term_pcp_cpu_jtag_debug_module AND pcp_cpu_jtag_debug_module_allgrants)) OR ((end_xfer_arb_share_counter_term_pcp_cpu_jtag_debug_module AND NOT pcp_cpu_jtag_debug_module_non_bursting_master_requests));
  --pcp_cpu_jtag_debug_module_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pcp_cpu_jtag_debug_module_arb_share_counter <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      if std_logic'(pcp_cpu_jtag_debug_module_arb_counter_enable) = '1' then 
        pcp_cpu_jtag_debug_module_arb_share_counter <= pcp_cpu_jtag_debug_module_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --pcp_cpu_jtag_debug_module_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pcp_cpu_jtag_debug_module_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((or_reduce(pcp_cpu_jtag_debug_module_master_qreq_vector) AND end_xfer_arb_share_counter_term_pcp_cpu_jtag_debug_module)) OR ((end_xfer_arb_share_counter_term_pcp_cpu_jtag_debug_module AND NOT pcp_cpu_jtag_debug_module_non_bursting_master_requests)))) = '1' then 
        pcp_cpu_jtag_debug_module_slavearbiterlockenable <= or_reduce(pcp_cpu_jtag_debug_module_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --pcp_cpu/data_master pcp_cpu/jtag_debug_module arbiterlock, which is an e_assign
  pcp_cpu_data_master_arbiterlock <= pcp_cpu_jtag_debug_module_slavearbiterlockenable AND pcp_cpu_data_master_continuerequest;
  --pcp_cpu_jtag_debug_module_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  pcp_cpu_jtag_debug_module_slavearbiterlockenable2 <= or_reduce(pcp_cpu_jtag_debug_module_arb_share_counter_next_value);
  --pcp_cpu/data_master pcp_cpu/jtag_debug_module arbiterlock2, which is an e_assign
  pcp_cpu_data_master_arbiterlock2 <= pcp_cpu_jtag_debug_module_slavearbiterlockenable2 AND pcp_cpu_data_master_continuerequest;
  --pcp_cpu/instruction_master pcp_cpu/jtag_debug_module arbiterlock, which is an e_assign
  pcp_cpu_instruction_master_arbiterlock <= pcp_cpu_jtag_debug_module_slavearbiterlockenable AND pcp_cpu_instruction_master_continuerequest;
  --pcp_cpu/instruction_master pcp_cpu/jtag_debug_module arbiterlock2, which is an e_assign
  pcp_cpu_instruction_master_arbiterlock2 <= pcp_cpu_jtag_debug_module_slavearbiterlockenable2 AND pcp_cpu_instruction_master_continuerequest;
  --pcp_cpu/instruction_master granted pcp_cpu/jtag_debug_module last time, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      last_cycle_pcp_cpu_instruction_master_granted_slave_pcp_cpu_jtag_debug_module <= std_logic'('0');
    elsif clk'event and clk = '1' then
      last_cycle_pcp_cpu_instruction_master_granted_slave_pcp_cpu_jtag_debug_module <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(pcp_cpu_instruction_master_saved_grant_pcp_cpu_jtag_debug_module) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((pcp_cpu_jtag_debug_module_arbitration_holdoff_internal OR NOT internal_pcp_cpu_instruction_master_requests_pcp_cpu_jtag_debug_module))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_pcp_cpu_instruction_master_granted_slave_pcp_cpu_jtag_debug_module))))));
    end if;

  end process;

  --pcp_cpu_instruction_master_continuerequest continued request, which is an e_mux
  pcp_cpu_instruction_master_continuerequest <= last_cycle_pcp_cpu_instruction_master_granted_slave_pcp_cpu_jtag_debug_module AND internal_pcp_cpu_instruction_master_requests_pcp_cpu_jtag_debug_module;
  --pcp_cpu_jtag_debug_module_any_continuerequest at least one master continues requesting, which is an e_mux
  pcp_cpu_jtag_debug_module_any_continuerequest <= pcp_cpu_instruction_master_continuerequest OR pcp_cpu_data_master_continuerequest;
  internal_pcp_cpu_data_master_qualified_request_pcp_cpu_jtag_debug_module <= internal_pcp_cpu_data_master_requests_pcp_cpu_jtag_debug_module AND NOT (((((NOT pcp_cpu_data_master_waitrequest) AND pcp_cpu_data_master_write)) OR pcp_cpu_instruction_master_arbiterlock));
  --pcp_cpu_jtag_debug_module_writedata mux, which is an e_mux
  pcp_cpu_jtag_debug_module_writedata <= pcp_cpu_data_master_writedata;
  internal_pcp_cpu_instruction_master_requests_pcp_cpu_jtag_debug_module <= ((to_std_logic(((Std_Logic_Vector'(pcp_cpu_instruction_master_address_to_slave(25 DOWNTO 11) & std_logic_vector'("00000000000")) = std_logic_vector'("00000000000001100000000000")))) AND (pcp_cpu_instruction_master_read))) AND pcp_cpu_instruction_master_read;
  --pcp_cpu/data_master granted pcp_cpu/jtag_debug_module last time, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      last_cycle_pcp_cpu_data_master_granted_slave_pcp_cpu_jtag_debug_module <= std_logic'('0');
    elsif clk'event and clk = '1' then
      last_cycle_pcp_cpu_data_master_granted_slave_pcp_cpu_jtag_debug_module <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(pcp_cpu_data_master_saved_grant_pcp_cpu_jtag_debug_module) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((pcp_cpu_jtag_debug_module_arbitration_holdoff_internal OR NOT internal_pcp_cpu_data_master_requests_pcp_cpu_jtag_debug_module))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_pcp_cpu_data_master_granted_slave_pcp_cpu_jtag_debug_module))))));
    end if;

  end process;

  --pcp_cpu_data_master_continuerequest continued request, which is an e_mux
  pcp_cpu_data_master_continuerequest <= last_cycle_pcp_cpu_data_master_granted_slave_pcp_cpu_jtag_debug_module AND internal_pcp_cpu_data_master_requests_pcp_cpu_jtag_debug_module;
  internal_pcp_cpu_instruction_master_qualified_request_pcp_cpu_jtag_debug_module <= internal_pcp_cpu_instruction_master_requests_pcp_cpu_jtag_debug_module AND NOT ((((pcp_cpu_instruction_master_read AND to_std_logic((((std_logic_vector'("000000000000000000000000000000") & (pcp_cpu_instruction_master_latency_counter)) /= std_logic_vector'("00000000000000000000000000000000")))))) OR pcp_cpu_data_master_arbiterlock));
  --local readdatavalid pcp_cpu_instruction_master_read_data_valid_pcp_cpu_jtag_debug_module, which is an e_mux
  pcp_cpu_instruction_master_read_data_valid_pcp_cpu_jtag_debug_module <= (internal_pcp_cpu_instruction_master_granted_pcp_cpu_jtag_debug_module AND pcp_cpu_instruction_master_read) AND NOT pcp_cpu_jtag_debug_module_waits_for_read;
  --allow new arb cycle for pcp_cpu/jtag_debug_module, which is an e_assign
  pcp_cpu_jtag_debug_module_allow_new_arb_cycle <= NOT pcp_cpu_data_master_arbiterlock AND NOT pcp_cpu_instruction_master_arbiterlock;
  --pcp_cpu/instruction_master assignment into master qualified-requests vector for pcp_cpu/jtag_debug_module, which is an e_assign
  pcp_cpu_jtag_debug_module_master_qreq_vector(0) <= internal_pcp_cpu_instruction_master_qualified_request_pcp_cpu_jtag_debug_module;
  --pcp_cpu/instruction_master grant pcp_cpu/jtag_debug_module, which is an e_assign
  internal_pcp_cpu_instruction_master_granted_pcp_cpu_jtag_debug_module <= pcp_cpu_jtag_debug_module_grant_vector(0);
  --pcp_cpu/instruction_master saved-grant pcp_cpu/jtag_debug_module, which is an e_assign
  pcp_cpu_instruction_master_saved_grant_pcp_cpu_jtag_debug_module <= pcp_cpu_jtag_debug_module_arb_winner(0) AND internal_pcp_cpu_instruction_master_requests_pcp_cpu_jtag_debug_module;
  --pcp_cpu/data_master assignment into master qualified-requests vector for pcp_cpu/jtag_debug_module, which is an e_assign
  pcp_cpu_jtag_debug_module_master_qreq_vector(1) <= internal_pcp_cpu_data_master_qualified_request_pcp_cpu_jtag_debug_module;
  --pcp_cpu/data_master grant pcp_cpu/jtag_debug_module, which is an e_assign
  internal_pcp_cpu_data_master_granted_pcp_cpu_jtag_debug_module <= pcp_cpu_jtag_debug_module_grant_vector(1);
  --pcp_cpu/data_master saved-grant pcp_cpu/jtag_debug_module, which is an e_assign
  pcp_cpu_data_master_saved_grant_pcp_cpu_jtag_debug_module <= pcp_cpu_jtag_debug_module_arb_winner(1) AND internal_pcp_cpu_data_master_requests_pcp_cpu_jtag_debug_module;
  --pcp_cpu/jtag_debug_module chosen-master double-vector, which is an e_assign
  pcp_cpu_jtag_debug_module_chosen_master_double_vector <= A_EXT (((std_logic_vector'("0") & ((pcp_cpu_jtag_debug_module_master_qreq_vector & pcp_cpu_jtag_debug_module_master_qreq_vector))) AND (((std_logic_vector'("0") & (Std_Logic_Vector'(NOT pcp_cpu_jtag_debug_module_master_qreq_vector & NOT pcp_cpu_jtag_debug_module_master_qreq_vector))) + (std_logic_vector'("000") & (pcp_cpu_jtag_debug_module_arb_addend))))), 4);
  --stable onehot encoding of arb winner
  pcp_cpu_jtag_debug_module_arb_winner <= A_WE_StdLogicVector((std_logic'(((pcp_cpu_jtag_debug_module_allow_new_arb_cycle AND or_reduce(pcp_cpu_jtag_debug_module_grant_vector)))) = '1'), pcp_cpu_jtag_debug_module_grant_vector, pcp_cpu_jtag_debug_module_saved_chosen_master_vector);
  --saved pcp_cpu_jtag_debug_module_grant_vector, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pcp_cpu_jtag_debug_module_saved_chosen_master_vector <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      if std_logic'(pcp_cpu_jtag_debug_module_allow_new_arb_cycle) = '1' then 
        pcp_cpu_jtag_debug_module_saved_chosen_master_vector <= A_WE_StdLogicVector((std_logic'(or_reduce(pcp_cpu_jtag_debug_module_grant_vector)) = '1'), pcp_cpu_jtag_debug_module_grant_vector, pcp_cpu_jtag_debug_module_saved_chosen_master_vector);
      end if;
    end if;

  end process;

  --onehot encoding of chosen master
  pcp_cpu_jtag_debug_module_grant_vector <= Std_Logic_Vector'(A_ToStdLogicVector(((pcp_cpu_jtag_debug_module_chosen_master_double_vector(1) OR pcp_cpu_jtag_debug_module_chosen_master_double_vector(3)))) & A_ToStdLogicVector(((pcp_cpu_jtag_debug_module_chosen_master_double_vector(0) OR pcp_cpu_jtag_debug_module_chosen_master_double_vector(2)))));
  --pcp_cpu/jtag_debug_module chosen master rotated left, which is an e_assign
  pcp_cpu_jtag_debug_module_chosen_master_rot_left <= A_EXT (A_WE_StdLogicVector((((A_SLL(pcp_cpu_jtag_debug_module_arb_winner,std_logic_vector'("00000000000000000000000000000001")))) /= std_logic_vector'("00")), (std_logic_vector'("000000000000000000000000000000") & ((A_SLL(pcp_cpu_jtag_debug_module_arb_winner,std_logic_vector'("00000000000000000000000000000001"))))), std_logic_vector'("00000000000000000000000000000001")), 2);
  --pcp_cpu/jtag_debug_module's addend for next-master-grant
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pcp_cpu_jtag_debug_module_arb_addend <= std_logic_vector'("01");
    elsif clk'event and clk = '1' then
      if std_logic'(or_reduce(pcp_cpu_jtag_debug_module_grant_vector)) = '1' then 
        pcp_cpu_jtag_debug_module_arb_addend <= A_WE_StdLogicVector((std_logic'(pcp_cpu_jtag_debug_module_end_xfer) = '1'), pcp_cpu_jtag_debug_module_chosen_master_rot_left, pcp_cpu_jtag_debug_module_grant_vector);
      end if;
    end if;

  end process;

  pcp_cpu_jtag_debug_module_begintransfer <= pcp_cpu_jtag_debug_module_begins_xfer;
  --pcp_cpu_jtag_debug_module_reset_n assignment, which is an e_assign
  pcp_cpu_jtag_debug_module_reset_n <= reset_n;
  --assign pcp_cpu_jtag_debug_module_resetrequest_from_sa = pcp_cpu_jtag_debug_module_resetrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  pcp_cpu_jtag_debug_module_resetrequest_from_sa <= pcp_cpu_jtag_debug_module_resetrequest;
  pcp_cpu_jtag_debug_module_chipselect <= internal_pcp_cpu_data_master_granted_pcp_cpu_jtag_debug_module OR internal_pcp_cpu_instruction_master_granted_pcp_cpu_jtag_debug_module;
  --pcp_cpu_jtag_debug_module_firsttransfer first transaction, which is an e_assign
  pcp_cpu_jtag_debug_module_firsttransfer <= A_WE_StdLogic((std_logic'(pcp_cpu_jtag_debug_module_begins_xfer) = '1'), pcp_cpu_jtag_debug_module_unreg_firsttransfer, pcp_cpu_jtag_debug_module_reg_firsttransfer);
  --pcp_cpu_jtag_debug_module_unreg_firsttransfer first transaction, which is an e_assign
  pcp_cpu_jtag_debug_module_unreg_firsttransfer <= NOT ((pcp_cpu_jtag_debug_module_slavearbiterlockenable AND pcp_cpu_jtag_debug_module_any_continuerequest));
  --pcp_cpu_jtag_debug_module_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pcp_cpu_jtag_debug_module_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(pcp_cpu_jtag_debug_module_begins_xfer) = '1' then 
        pcp_cpu_jtag_debug_module_reg_firsttransfer <= pcp_cpu_jtag_debug_module_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --pcp_cpu_jtag_debug_module_beginbursttransfer_internal begin burst transfer, which is an e_assign
  pcp_cpu_jtag_debug_module_beginbursttransfer_internal <= pcp_cpu_jtag_debug_module_begins_xfer;
  --pcp_cpu_jtag_debug_module_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  pcp_cpu_jtag_debug_module_arbitration_holdoff_internal <= pcp_cpu_jtag_debug_module_begins_xfer AND pcp_cpu_jtag_debug_module_firsttransfer;
  --pcp_cpu_jtag_debug_module_write assignment, which is an e_mux
  pcp_cpu_jtag_debug_module_write <= internal_pcp_cpu_data_master_granted_pcp_cpu_jtag_debug_module AND pcp_cpu_data_master_write;
  shifted_address_to_pcp_cpu_jtag_debug_module_from_pcp_cpu_data_master <= pcp_cpu_data_master_address_to_slave;
  --pcp_cpu_jtag_debug_module_address mux, which is an e_mux
  pcp_cpu_jtag_debug_module_address <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_pcp_cpu_data_master_granted_pcp_cpu_jtag_debug_module)) = '1'), (A_SRL(shifted_address_to_pcp_cpu_jtag_debug_module_from_pcp_cpu_data_master,std_logic_vector'("00000000000000000000000000000010"))), (A_SRL(shifted_address_to_pcp_cpu_jtag_debug_module_from_pcp_cpu_instruction_master,std_logic_vector'("00000000000000000000000000000010")))), 9);
  shifted_address_to_pcp_cpu_jtag_debug_module_from_pcp_cpu_instruction_master <= pcp_cpu_instruction_master_address_to_slave;
  --d1_pcp_cpu_jtag_debug_module_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_pcp_cpu_jtag_debug_module_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_pcp_cpu_jtag_debug_module_end_xfer <= pcp_cpu_jtag_debug_module_end_xfer;
    end if;

  end process;

  --pcp_cpu_jtag_debug_module_waits_for_read in a cycle, which is an e_mux
  pcp_cpu_jtag_debug_module_waits_for_read <= pcp_cpu_jtag_debug_module_in_a_read_cycle AND pcp_cpu_jtag_debug_module_begins_xfer;
  --pcp_cpu_jtag_debug_module_in_a_read_cycle assignment, which is an e_assign
  pcp_cpu_jtag_debug_module_in_a_read_cycle <= ((internal_pcp_cpu_data_master_granted_pcp_cpu_jtag_debug_module AND pcp_cpu_data_master_read)) OR ((internal_pcp_cpu_instruction_master_granted_pcp_cpu_jtag_debug_module AND pcp_cpu_instruction_master_read));
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= pcp_cpu_jtag_debug_module_in_a_read_cycle;
  --pcp_cpu_jtag_debug_module_waits_for_write in a cycle, which is an e_mux
  pcp_cpu_jtag_debug_module_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pcp_cpu_jtag_debug_module_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --pcp_cpu_jtag_debug_module_in_a_write_cycle assignment, which is an e_assign
  pcp_cpu_jtag_debug_module_in_a_write_cycle <= internal_pcp_cpu_data_master_granted_pcp_cpu_jtag_debug_module AND pcp_cpu_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= pcp_cpu_jtag_debug_module_in_a_write_cycle;
  wait_for_pcp_cpu_jtag_debug_module_counter <= std_logic'('0');
  --pcp_cpu_jtag_debug_module_byteenable byte enable port mux, which is an e_mux
  pcp_cpu_jtag_debug_module_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_pcp_cpu_data_master_granted_pcp_cpu_jtag_debug_module)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (pcp_cpu_data_master_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))), 4);
  --debugaccess mux, which is an e_mux
  pcp_cpu_jtag_debug_module_debugaccess <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((internal_pcp_cpu_data_master_granted_pcp_cpu_jtag_debug_module)) = '1'), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pcp_cpu_data_master_debugaccess))), std_logic_vector'("00000000000000000000000000000000")));
  --vhdl renameroo for output signals
  pcp_cpu_data_master_granted_pcp_cpu_jtag_debug_module <= internal_pcp_cpu_data_master_granted_pcp_cpu_jtag_debug_module;
  --vhdl renameroo for output signals
  pcp_cpu_data_master_qualified_request_pcp_cpu_jtag_debug_module <= internal_pcp_cpu_data_master_qualified_request_pcp_cpu_jtag_debug_module;
  --vhdl renameroo for output signals
  pcp_cpu_data_master_requests_pcp_cpu_jtag_debug_module <= internal_pcp_cpu_data_master_requests_pcp_cpu_jtag_debug_module;
  --vhdl renameroo for output signals
  pcp_cpu_instruction_master_granted_pcp_cpu_jtag_debug_module <= internal_pcp_cpu_instruction_master_granted_pcp_cpu_jtag_debug_module;
  --vhdl renameroo for output signals
  pcp_cpu_instruction_master_qualified_request_pcp_cpu_jtag_debug_module <= internal_pcp_cpu_instruction_master_qualified_request_pcp_cpu_jtag_debug_module;
  --vhdl renameroo for output signals
  pcp_cpu_instruction_master_requests_pcp_cpu_jtag_debug_module <= internal_pcp_cpu_instruction_master_requests_pcp_cpu_jtag_debug_module;
--synthesis translate_off
    --pcp_cpu/jtag_debug_module enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --grant signals are active simultaneously, which is an e_process
    process (clk)
    VARIABLE write_line43 : line;
    begin
      if clk'event and clk = '1' then
        if (std_logic_vector'("000000000000000000000000000000") & (((std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(internal_pcp_cpu_data_master_granted_pcp_cpu_jtag_debug_module))) + (std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(internal_pcp_cpu_instruction_master_granted_pcp_cpu_jtag_debug_module))))))>std_logic_vector'("00000000000000000000000000000001") then 
          write(write_line43, now);
          write(write_line43, string'(": "));
          write(write_line43, string'("> 1 of grant signals are active simultaneously"));
          write(output, write_line43.all);
          deallocate (write_line43);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --saved_grant signals are active simultaneously, which is an e_process
    process (clk)
    VARIABLE write_line44 : line;
    begin
      if clk'event and clk = '1' then
        if (std_logic_vector'("000000000000000000000000000000") & (((std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(pcp_cpu_data_master_saved_grant_pcp_cpu_jtag_debug_module))) + (std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(pcp_cpu_instruction_master_saved_grant_pcp_cpu_jtag_debug_module))))))>std_logic_vector'("00000000000000000000000000000001") then 
          write(write_line44, now);
          write(write_line44, string'(": "));
          write(write_line44, string'("> 1 of saved_grant signals are active simultaneously"));
          write(output, write_line44.all);
          deallocate (write_line44);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity OpenMAC_0_CMP_irq_from_sa_clock_crossing_pcp_cpu_data_master_module is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC
              );
end entity OpenMAC_0_CMP_irq_from_sa_clock_crossing_pcp_cpu_data_master_module;


architecture europa of OpenMAC_0_CMP_irq_from_sa_clock_crossing_pcp_cpu_data_master_module is
                signal data_in_d1 :  STD_LOGIC;
attribute ALTERA_ATTRIBUTE : string;
attribute ALTERA_ATTRIBUTE of data_in_d1 : signal is "{-from ""*""} CUT=ON ; PRESERVE_REGISTER=ON";
attribute ALTERA_ATTRIBUTE of data_out : signal is "PRESERVE_REGISTER=ON";

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      data_in_d1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      data_in_d1 <= data_in;
    end if;

  end process;

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      data_out <= std_logic'('0');
    elsif clk'event and clk = '1' then
      data_out <= data_in_d1;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity OpenMAC_0_REG_irq_from_sa_clock_crossing_pcp_cpu_data_master_module is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC
              );
end entity OpenMAC_0_REG_irq_from_sa_clock_crossing_pcp_cpu_data_master_module;


architecture europa of OpenMAC_0_REG_irq_from_sa_clock_crossing_pcp_cpu_data_master_module is
                signal data_in_d1 :  STD_LOGIC;
attribute ALTERA_ATTRIBUTE : string;
attribute ALTERA_ATTRIBUTE of data_in_d1 : signal is "{-from ""*""} CUT=ON ; PRESERVE_REGISTER=ON";
attribute ALTERA_ATTRIBUTE of data_out : signal is "PRESERVE_REGISTER=ON";

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      data_in_d1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      data_in_d1 <= data_in;
    end if;

  end process;

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      data_out <= std_logic'('0');
    elsif clk'event and clk = '1' then
      data_out <= data_in_d1;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity jtag_uart_0_avalon_jtag_slave_irq_from_sa_clock_crossing_pcp_cpu_data_master_module is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC
              );
end entity jtag_uart_0_avalon_jtag_slave_irq_from_sa_clock_crossing_pcp_cpu_data_master_module;


architecture europa of jtag_uart_0_avalon_jtag_slave_irq_from_sa_clock_crossing_pcp_cpu_data_master_module is
                signal data_in_d1 :  STD_LOGIC;
attribute ALTERA_ATTRIBUTE : string;
attribute ALTERA_ATTRIBUTE of data_in_d1 : signal is "{-from ""*""} CUT=ON ; PRESERVE_REGISTER=ON";
attribute ALTERA_ATTRIBUTE of data_out : signal is "PRESERVE_REGISTER=ON";

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      data_in_d1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      data_in_d1 <= data_in;
    end if;

  end process;

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      data_out <= std_logic'('0');
    elsif clk'event and clk = '1' then
      data_out <= data_in_d1;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity system_timer_s1_irq_from_sa_clock_crossing_pcp_cpu_data_master_module is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC
              );
end entity system_timer_s1_irq_from_sa_clock_crossing_pcp_cpu_data_master_module;


architecture europa of system_timer_s1_irq_from_sa_clock_crossing_pcp_cpu_data_master_module is
                signal data_in_d1 :  STD_LOGIC;
attribute ALTERA_ATTRIBUTE : string;
attribute ALTERA_ATTRIBUTE of data_in_d1 : signal is "{-from ""*""} CUT=ON ; PRESERVE_REGISTER=ON";
attribute ALTERA_ATTRIBUTE of data_out : signal is "PRESERVE_REGISTER=ON";

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      data_in_d1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      data_in_d1 <= data_in;
    end if;

  end process;

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      data_out <= std_logic'('0');
    elsif clk'event and clk = '1' then
      data_out <= data_in_d1;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity pcp_cpu_data_master_arbitrator is 
        port (
              -- inputs:
                 signal DBC3C40_SRAM_0_avalon_tristate_slave_wait_counter_eq_0 : IN STD_LOGIC;
                 signal OpenMAC_0_CMP_irq_from_sa : IN STD_LOGIC;
                 signal OpenMAC_0_REG_irq_from_sa : IN STD_LOGIC;
                 signal OpenMAC_0_iBuf_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal OpenMAC_0_iBuf_wait_counter_eq_0 : IN STD_LOGIC;
                 signal cfi_flash_0_s1_wait_counter_eq_0 : IN STD_LOGIC;
                 signal cfi_flash_0_s1_wait_counter_eq_1 : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal clk90Meg : IN STD_LOGIC;
                 signal clk90Meg_reset_n : IN STD_LOGIC;
                 signal clock_crossing_0_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal clock_crossing_0_s1_waitrequest_from_sa : IN STD_LOGIC;
                 signal cnApi_Av2Av_0_pcp_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal cnApi_Av2Av_0_pcp_wait_counter_eq_0 : IN STD_LOGIC;
                 signal d1_OpenMAC_0_iBuf_end_xfer : IN STD_LOGIC;
                 signal d1_clock_crossing_0_s1_end_xfer : IN STD_LOGIC;
                 signal d1_cnApi_Av2Av_0_pcp_end_xfer : IN STD_LOGIC;
                 signal d1_epcs_flash_controller_0_epcs_control_port_end_xfer : IN STD_LOGIC;
                 signal d1_niosII_openMac_clock_0_in_end_xfer : IN STD_LOGIC;
                 signal d1_niosII_openMac_clock_1_in_end_xfer : IN STD_LOGIC;
                 signal d1_niosII_openMac_clock_2_in_end_xfer : IN STD_LOGIC;
                 signal d1_niosII_openMac_clock_3_in_end_xfer : IN STD_LOGIC;
                 signal d1_niosII_openMac_clock_4_in_end_xfer : IN STD_LOGIC;
                 signal d1_onchip_memory_0_s1_end_xfer : IN STD_LOGIC;
                 signal d1_pcp_cpu_jtag_debug_module_end_xfer : IN STD_LOGIC;
                 signal d1_tri_state_bridge_0_avalon_slave_end_xfer : IN STD_LOGIC;
                 signal epcs_flash_controller_0_epcs_control_port_irq_from_sa : IN STD_LOGIC;
                 signal epcs_flash_controller_0_epcs_control_port_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal incoming_tri_state_bridge_0_data : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal incoming_tri_state_bridge_0_data_with_Xs_converted_to_0 : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal jtag_uart_0_avalon_jtag_slave_irq_from_sa : IN STD_LOGIC;
                 signal niosII_openMac_clock_0_in_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal niosII_openMac_clock_0_in_waitrequest_from_sa : IN STD_LOGIC;
                 signal niosII_openMac_clock_1_in_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal niosII_openMac_clock_1_in_waitrequest_from_sa : IN STD_LOGIC;
                 signal niosII_openMac_clock_2_in_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal niosII_openMac_clock_2_in_waitrequest_from_sa : IN STD_LOGIC;
                 signal niosII_openMac_clock_3_in_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal niosII_openMac_clock_3_in_waitrequest_from_sa : IN STD_LOGIC;
                 signal niosII_openMac_clock_4_in_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal niosII_openMac_clock_4_in_waitrequest_from_sa : IN STD_LOGIC;
                 signal onchip_memory_0_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal pcp_cpu_data_master_address : IN STD_LOGIC_VECTOR (25 DOWNTO 0);
                 signal pcp_cpu_data_master_byteenable_DBC3C40_SRAM_0_avalon_tristate_slave : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal pcp_cpu_data_master_byteenable_cfi_flash_0_s1 : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal pcp_cpu_data_master_byteenable_niosII_openMac_clock_2_in : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal pcp_cpu_data_master_granted_DBC3C40_SRAM_0_avalon_tristate_slave : IN STD_LOGIC;
                 signal pcp_cpu_data_master_granted_OpenMAC_0_iBuf : IN STD_LOGIC;
                 signal pcp_cpu_data_master_granted_cfi_flash_0_s1 : IN STD_LOGIC;
                 signal pcp_cpu_data_master_granted_clock_crossing_0_s1 : IN STD_LOGIC;
                 signal pcp_cpu_data_master_granted_cnApi_Av2Av_0_pcp : IN STD_LOGIC;
                 signal pcp_cpu_data_master_granted_epcs_flash_controller_0_epcs_control_port : IN STD_LOGIC;
                 signal pcp_cpu_data_master_granted_niosII_openMac_clock_0_in : IN STD_LOGIC;
                 signal pcp_cpu_data_master_granted_niosII_openMac_clock_1_in : IN STD_LOGIC;
                 signal pcp_cpu_data_master_granted_niosII_openMac_clock_2_in : IN STD_LOGIC;
                 signal pcp_cpu_data_master_granted_niosII_openMac_clock_3_in : IN STD_LOGIC;
                 signal pcp_cpu_data_master_granted_niosII_openMac_clock_4_in : IN STD_LOGIC;
                 signal pcp_cpu_data_master_granted_onchip_memory_0_s1 : IN STD_LOGIC;
                 signal pcp_cpu_data_master_granted_pcp_cpu_jtag_debug_module : IN STD_LOGIC;
                 signal pcp_cpu_data_master_qualified_request_DBC3C40_SRAM_0_avalon_tristate_slave : IN STD_LOGIC;
                 signal pcp_cpu_data_master_qualified_request_OpenMAC_0_iBuf : IN STD_LOGIC;
                 signal pcp_cpu_data_master_qualified_request_cfi_flash_0_s1 : IN STD_LOGIC;
                 signal pcp_cpu_data_master_qualified_request_clock_crossing_0_s1 : IN STD_LOGIC;
                 signal pcp_cpu_data_master_qualified_request_cnApi_Av2Av_0_pcp : IN STD_LOGIC;
                 signal pcp_cpu_data_master_qualified_request_epcs_flash_controller_0_epcs_control_port : IN STD_LOGIC;
                 signal pcp_cpu_data_master_qualified_request_niosII_openMac_clock_0_in : IN STD_LOGIC;
                 signal pcp_cpu_data_master_qualified_request_niosII_openMac_clock_1_in : IN STD_LOGIC;
                 signal pcp_cpu_data_master_qualified_request_niosII_openMac_clock_2_in : IN STD_LOGIC;
                 signal pcp_cpu_data_master_qualified_request_niosII_openMac_clock_3_in : IN STD_LOGIC;
                 signal pcp_cpu_data_master_qualified_request_niosII_openMac_clock_4_in : IN STD_LOGIC;
                 signal pcp_cpu_data_master_qualified_request_onchip_memory_0_s1 : IN STD_LOGIC;
                 signal pcp_cpu_data_master_qualified_request_pcp_cpu_jtag_debug_module : IN STD_LOGIC;
                 signal pcp_cpu_data_master_read : IN STD_LOGIC;
                 signal pcp_cpu_data_master_read_data_valid_DBC3C40_SRAM_0_avalon_tristate_slave : IN STD_LOGIC;
                 signal pcp_cpu_data_master_read_data_valid_OpenMAC_0_iBuf : IN STD_LOGIC;
                 signal pcp_cpu_data_master_read_data_valid_cfi_flash_0_s1 : IN STD_LOGIC;
                 signal pcp_cpu_data_master_read_data_valid_clock_crossing_0_s1 : IN STD_LOGIC;
                 signal pcp_cpu_data_master_read_data_valid_clock_crossing_0_s1_shift_register : IN STD_LOGIC;
                 signal pcp_cpu_data_master_read_data_valid_cnApi_Av2Av_0_pcp : IN STD_LOGIC;
                 signal pcp_cpu_data_master_read_data_valid_epcs_flash_controller_0_epcs_control_port : IN STD_LOGIC;
                 signal pcp_cpu_data_master_read_data_valid_niosII_openMac_clock_0_in : IN STD_LOGIC;
                 signal pcp_cpu_data_master_read_data_valid_niosII_openMac_clock_1_in : IN STD_LOGIC;
                 signal pcp_cpu_data_master_read_data_valid_niosII_openMac_clock_2_in : IN STD_LOGIC;
                 signal pcp_cpu_data_master_read_data_valid_niosII_openMac_clock_3_in : IN STD_LOGIC;
                 signal pcp_cpu_data_master_read_data_valid_niosII_openMac_clock_4_in : IN STD_LOGIC;
                 signal pcp_cpu_data_master_read_data_valid_onchip_memory_0_s1 : IN STD_LOGIC;
                 signal pcp_cpu_data_master_read_data_valid_pcp_cpu_jtag_debug_module : IN STD_LOGIC;
                 signal pcp_cpu_data_master_requests_DBC3C40_SRAM_0_avalon_tristate_slave : IN STD_LOGIC;
                 signal pcp_cpu_data_master_requests_OpenMAC_0_iBuf : IN STD_LOGIC;
                 signal pcp_cpu_data_master_requests_cfi_flash_0_s1 : IN STD_LOGIC;
                 signal pcp_cpu_data_master_requests_clock_crossing_0_s1 : IN STD_LOGIC;
                 signal pcp_cpu_data_master_requests_cnApi_Av2Av_0_pcp : IN STD_LOGIC;
                 signal pcp_cpu_data_master_requests_epcs_flash_controller_0_epcs_control_port : IN STD_LOGIC;
                 signal pcp_cpu_data_master_requests_niosII_openMac_clock_0_in : IN STD_LOGIC;
                 signal pcp_cpu_data_master_requests_niosII_openMac_clock_1_in : IN STD_LOGIC;
                 signal pcp_cpu_data_master_requests_niosII_openMac_clock_2_in : IN STD_LOGIC;
                 signal pcp_cpu_data_master_requests_niosII_openMac_clock_3_in : IN STD_LOGIC;
                 signal pcp_cpu_data_master_requests_niosII_openMac_clock_4_in : IN STD_LOGIC;
                 signal pcp_cpu_data_master_requests_onchip_memory_0_s1 : IN STD_LOGIC;
                 signal pcp_cpu_data_master_requests_pcp_cpu_jtag_debug_module : IN STD_LOGIC;
                 signal pcp_cpu_data_master_write : IN STD_LOGIC;
                 signal pcp_cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal pcp_cpu_jtag_debug_module_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal registered_pcp_cpu_data_master_read_data_valid_DBC3C40_SRAM_0_avalon_tristate_slave : IN STD_LOGIC;
                 signal registered_pcp_cpu_data_master_read_data_valid_cfi_flash_0_s1 : IN STD_LOGIC;
                 signal registered_pcp_cpu_data_master_read_data_valid_onchip_memory_0_s1 : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal system_timer_s1_irq_from_sa : IN STD_LOGIC;

              -- outputs:
                 signal pcp_cpu_data_master_address_to_slave : OUT STD_LOGIC_VECTOR (25 DOWNTO 0);
                 signal pcp_cpu_data_master_dbs_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal pcp_cpu_data_master_dbs_write_16 : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal pcp_cpu_data_master_irq : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal pcp_cpu_data_master_no_byte_enables_and_last_term : OUT STD_LOGIC;
                 signal pcp_cpu_data_master_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal pcp_cpu_data_master_waitrequest : OUT STD_LOGIC
              );
end entity pcp_cpu_data_master_arbitrator;


architecture europa of pcp_cpu_data_master_arbitrator is
component OpenMAC_0_CMP_irq_from_sa_clock_crossing_pcp_cpu_data_master_module is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC
                 );
end component OpenMAC_0_CMP_irq_from_sa_clock_crossing_pcp_cpu_data_master_module;

component OpenMAC_0_REG_irq_from_sa_clock_crossing_pcp_cpu_data_master_module is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC
                 );
end component OpenMAC_0_REG_irq_from_sa_clock_crossing_pcp_cpu_data_master_module;

component jtag_uart_0_avalon_jtag_slave_irq_from_sa_clock_crossing_pcp_cpu_data_master_module is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC
                 );
end component jtag_uart_0_avalon_jtag_slave_irq_from_sa_clock_crossing_pcp_cpu_data_master_module;

component system_timer_s1_irq_from_sa_clock_crossing_pcp_cpu_data_master_module is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC
                 );
end component system_timer_s1_irq_from_sa_clock_crossing_pcp_cpu_data_master_module;

                signal clk90Meg_OpenMAC_0_CMP_irq_from_sa :  STD_LOGIC;
                signal clk90Meg_OpenMAC_0_REG_irq_from_sa :  STD_LOGIC;
                signal clk90Meg_jtag_uart_0_avalon_jtag_slave_irq_from_sa :  STD_LOGIC;
                signal clk90Meg_system_timer_s1_irq_from_sa :  STD_LOGIC;
                signal dbs_16_reg_segment_0 :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal dbs_count_enable :  STD_LOGIC;
                signal dbs_counter_overflow :  STD_LOGIC;
                signal internal_pcp_cpu_data_master_address_to_slave :  STD_LOGIC_VECTOR (25 DOWNTO 0);
                signal internal_pcp_cpu_data_master_dbs_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal internal_pcp_cpu_data_master_no_byte_enables_and_last_term :  STD_LOGIC;
                signal internal_pcp_cpu_data_master_waitrequest :  STD_LOGIC;
                signal last_dbs_term_and_run :  STD_LOGIC;
                signal next_dbs_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal p1_dbs_16_reg_segment_0 :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal p1_registered_pcp_cpu_data_master_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal pcp_cpu_data_master_dbs_increment :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal pcp_cpu_data_master_run :  STD_LOGIC;
                signal pre_dbs_count_enable :  STD_LOGIC;
                signal r_0 :  STD_LOGIC;
                signal r_1 :  STD_LOGIC;
                signal r_2 :  STD_LOGIC;
                signal registered_pcp_cpu_data_master_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);

begin

  --r_0 master_run cascaded wait assignment, which is an e_assign
  r_0 <= Vector_To_Std_Logic((((((((((((((((((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pcp_cpu_data_master_qualified_request_OpenMAC_0_iBuf OR NOT pcp_cpu_data_master_requests_OpenMAC_0_iBuf)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT pcp_cpu_data_master_qualified_request_OpenMAC_0_iBuf OR NOT pcp_cpu_data_master_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT d1_OpenMAC_0_iBuf_end_xfer)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pcp_cpu_data_master_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT pcp_cpu_data_master_qualified_request_OpenMAC_0_iBuf OR NOT pcp_cpu_data_master_write)))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pcp_cpu_data_master_write)))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((pcp_cpu_data_master_qualified_request_clock_crossing_0_s1 OR pcp_cpu_data_master_read_data_valid_clock_crossing_0_s1) OR NOT pcp_cpu_data_master_requests_clock_crossing_0_s1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((NOT pcp_cpu_data_master_qualified_request_clock_crossing_0_s1 OR NOT pcp_cpu_data_master_read) OR ((pcp_cpu_data_master_read_data_valid_clock_crossing_0_s1 AND pcp_cpu_data_master_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT pcp_cpu_data_master_qualified_request_clock_crossing_0_s1 OR NOT ((pcp_cpu_data_master_read OR pcp_cpu_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT clock_crossing_0_s1_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pcp_cpu_data_master_read OR pcp_cpu_data_master_write)))))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pcp_cpu_data_master_qualified_request_cnApi_Av2Av_0_pcp OR NOT pcp_cpu_data_master_requests_cnApi_Av2Av_0_pcp)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT pcp_cpu_data_master_qualified_request_cnApi_Av2Av_0_pcp OR NOT pcp_cpu_data_master_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT d1_cnApi_Av2Av_0_pcp_end_xfer)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pcp_cpu_data_master_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT pcp_cpu_data_master_qualified_request_cnApi_Av2Av_0_pcp OR NOT pcp_cpu_data_master_write)))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pcp_cpu_data_master_write)))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pcp_cpu_data_master_qualified_request_epcs_flash_controller_0_epcs_control_port OR NOT pcp_cpu_data_master_requests_epcs_flash_controller_0_epcs_control_port)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pcp_cpu_data_master_granted_epcs_flash_controller_0_epcs_control_port OR NOT pcp_cpu_data_master_qualified_request_epcs_flash_controller_0_epcs_control_port)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT pcp_cpu_data_master_qualified_request_epcs_flash_controller_0_epcs_control_port OR NOT ((pcp_cpu_data_master_read OR pcp_cpu_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pcp_cpu_data_master_read OR pcp_cpu_data_master_write)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT pcp_cpu_data_master_qualified_request_epcs_flash_controller_0_epcs_control_port OR NOT ((pcp_cpu_data_master_read OR pcp_cpu_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pcp_cpu_data_master_read OR pcp_cpu_data_master_write)))))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pcp_cpu_data_master_qualified_request_niosII_openMac_clock_0_in OR NOT pcp_cpu_data_master_requests_niosII_openMac_clock_0_in)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT pcp_cpu_data_master_qualified_request_niosII_openMac_clock_0_in OR NOT ((pcp_cpu_data_master_read OR pcp_cpu_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT niosII_openMac_clock_0_in_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pcp_cpu_data_master_read OR pcp_cpu_data_master_write)))))))))));
  --cascaded wait assignment, which is an e_assign
  pcp_cpu_data_master_run <= (r_0 AND r_1) AND r_2;
  --r_1 master_run cascaded wait assignment, which is an e_assign
  r_1 <= Vector_To_Std_Logic(((((((((((((((((((((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT pcp_cpu_data_master_qualified_request_niosII_openMac_clock_0_in OR NOT ((pcp_cpu_data_master_read OR pcp_cpu_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT niosII_openMac_clock_0_in_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pcp_cpu_data_master_read OR pcp_cpu_data_master_write))))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pcp_cpu_data_master_qualified_request_niosII_openMac_clock_1_in OR NOT pcp_cpu_data_master_requests_niosII_openMac_clock_1_in)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT pcp_cpu_data_master_qualified_request_niosII_openMac_clock_1_in OR NOT ((pcp_cpu_data_master_read OR pcp_cpu_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT niosII_openMac_clock_1_in_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pcp_cpu_data_master_read OR pcp_cpu_data_master_write)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT pcp_cpu_data_master_qualified_request_niosII_openMac_clock_1_in OR NOT ((pcp_cpu_data_master_read OR pcp_cpu_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT niosII_openMac_clock_1_in_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pcp_cpu_data_master_read OR pcp_cpu_data_master_write)))))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((pcp_cpu_data_master_qualified_request_niosII_openMac_clock_2_in OR (((pcp_cpu_data_master_write AND NOT(or_reduce(pcp_cpu_data_master_byteenable_niosII_openMac_clock_2_in))) AND internal_pcp_cpu_data_master_dbs_address(1)))) OR NOT pcp_cpu_data_master_requests_niosII_openMac_clock_2_in)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT pcp_cpu_data_master_qualified_request_niosII_openMac_clock_2_in OR NOT pcp_cpu_data_master_read)))) OR ((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT niosII_openMac_clock_2_in_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((internal_pcp_cpu_data_master_dbs_address(1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pcp_cpu_data_master_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT pcp_cpu_data_master_qualified_request_niosII_openMac_clock_2_in OR NOT pcp_cpu_data_master_write)))) OR ((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT niosII_openMac_clock_2_in_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((internal_pcp_cpu_data_master_dbs_address(1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pcp_cpu_data_master_write)))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pcp_cpu_data_master_qualified_request_niosII_openMac_clock_3_in OR NOT pcp_cpu_data_master_requests_niosII_openMac_clock_3_in)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT pcp_cpu_data_master_qualified_request_niosII_openMac_clock_3_in OR NOT ((pcp_cpu_data_master_read OR pcp_cpu_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT niosII_openMac_clock_3_in_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pcp_cpu_data_master_read OR pcp_cpu_data_master_write)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT pcp_cpu_data_master_qualified_request_niosII_openMac_clock_3_in OR NOT ((pcp_cpu_data_master_read OR pcp_cpu_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT niosII_openMac_clock_3_in_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pcp_cpu_data_master_read OR pcp_cpu_data_master_write)))))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pcp_cpu_data_master_qualified_request_niosII_openMac_clock_4_in OR NOT pcp_cpu_data_master_requests_niosII_openMac_clock_4_in)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT pcp_cpu_data_master_qualified_request_niosII_openMac_clock_4_in OR NOT ((pcp_cpu_data_master_read OR pcp_cpu_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT niosII_openMac_clock_4_in_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pcp_cpu_data_master_read OR pcp_cpu_data_master_write)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT pcp_cpu_data_master_qualified_request_niosII_openMac_clock_4_in OR NOT ((pcp_cpu_data_master_read OR pcp_cpu_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT niosII_openMac_clock_4_in_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pcp_cpu_data_master_read OR pcp_cpu_data_master_write)))))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((pcp_cpu_data_master_qualified_request_onchip_memory_0_s1 OR registered_pcp_cpu_data_master_read_data_valid_onchip_memory_0_s1) OR NOT pcp_cpu_data_master_requests_onchip_memory_0_s1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pcp_cpu_data_master_granted_onchip_memory_0_s1 OR NOT pcp_cpu_data_master_qualified_request_onchip_memory_0_s1)))))));
  --r_2 master_run cascaded wait assignment, which is an e_assign
  r_2 <= Vector_To_Std_Logic(((((((((((((((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((NOT pcp_cpu_data_master_qualified_request_onchip_memory_0_s1 OR NOT pcp_cpu_data_master_read) OR ((registered_pcp_cpu_data_master_read_data_valid_onchip_memory_0_s1 AND pcp_cpu_data_master_read))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT pcp_cpu_data_master_qualified_request_onchip_memory_0_s1 OR NOT ((pcp_cpu_data_master_read OR pcp_cpu_data_master_write)))))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pcp_cpu_data_master_read OR pcp_cpu_data_master_write)))))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pcp_cpu_data_master_qualified_request_pcp_cpu_jtag_debug_module OR NOT pcp_cpu_data_master_requests_pcp_cpu_jtag_debug_module)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pcp_cpu_data_master_granted_pcp_cpu_jtag_debug_module OR NOT pcp_cpu_data_master_qualified_request_pcp_cpu_jtag_debug_module)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT pcp_cpu_data_master_qualified_request_pcp_cpu_jtag_debug_module OR NOT pcp_cpu_data_master_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pcp_cpu_data_master_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT pcp_cpu_data_master_qualified_request_pcp_cpu_jtag_debug_module OR NOT pcp_cpu_data_master_write)))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pcp_cpu_data_master_write)))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((((pcp_cpu_data_master_qualified_request_DBC3C40_SRAM_0_avalon_tristate_slave OR ((registered_pcp_cpu_data_master_read_data_valid_DBC3C40_SRAM_0_avalon_tristate_slave AND internal_pcp_cpu_data_master_dbs_address(1)))) OR (((pcp_cpu_data_master_write AND NOT(or_reduce(pcp_cpu_data_master_byteenable_DBC3C40_SRAM_0_avalon_tristate_slave))) AND internal_pcp_cpu_data_master_dbs_address(1)))) OR NOT pcp_cpu_data_master_requests_DBC3C40_SRAM_0_avalon_tristate_slave)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((((pcp_cpu_data_master_qualified_request_cfi_flash_0_s1 OR ((registered_pcp_cpu_data_master_read_data_valid_cfi_flash_0_s1 AND internal_pcp_cpu_data_master_dbs_address(1)))) OR (((pcp_cpu_data_master_write AND NOT(or_reduce(pcp_cpu_data_master_byteenable_cfi_flash_0_s1))) AND internal_pcp_cpu_data_master_dbs_address(1)))) OR NOT pcp_cpu_data_master_requests_cfi_flash_0_s1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pcp_cpu_data_master_granted_DBC3C40_SRAM_0_avalon_tristate_slave OR NOT pcp_cpu_data_master_qualified_request_DBC3C40_SRAM_0_avalon_tristate_slave)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pcp_cpu_data_master_granted_cfi_flash_0_s1 OR NOT pcp_cpu_data_master_qualified_request_cfi_flash_0_s1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((NOT pcp_cpu_data_master_qualified_request_DBC3C40_SRAM_0_avalon_tristate_slave OR NOT pcp_cpu_data_master_read) OR (((registered_pcp_cpu_data_master_read_data_valid_DBC3C40_SRAM_0_avalon_tristate_slave AND (internal_pcp_cpu_data_master_dbs_address(1))) AND pcp_cpu_data_master_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT pcp_cpu_data_master_qualified_request_DBC3C40_SRAM_0_avalon_tristate_slave OR NOT pcp_cpu_data_master_write)))) OR ((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT d1_tri_state_bridge_0_avalon_slave_end_xfer)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((internal_pcp_cpu_data_master_dbs_address(1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pcp_cpu_data_master_write)))))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((NOT pcp_cpu_data_master_qualified_request_cfi_flash_0_s1 OR NOT pcp_cpu_data_master_read) OR (((registered_pcp_cpu_data_master_read_data_valid_cfi_flash_0_s1 AND (internal_pcp_cpu_data_master_dbs_address(1))) AND pcp_cpu_data_master_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT pcp_cpu_data_master_qualified_request_cfi_flash_0_s1 OR NOT pcp_cpu_data_master_write)))) OR ((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cfi_flash_0_s1_wait_counter_eq_1)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((internal_pcp_cpu_data_master_dbs_address(1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pcp_cpu_data_master_write)))))))));
  --OpenMAC_0_CMP_irq_from_sa from clk50Meg to clk90Meg
  OpenMAC_0_CMP_irq_from_sa_clock_crossing_pcp_cpu_data_master : OpenMAC_0_CMP_irq_from_sa_clock_crossing_pcp_cpu_data_master_module
    port map(
      data_out => clk90Meg_OpenMAC_0_CMP_irq_from_sa,
      clk => clk90Meg,
      data_in => OpenMAC_0_CMP_irq_from_sa,
      reset_n => clk90Meg_reset_n
    );


  --irq assign, which is an e_assign
  pcp_cpu_data_master_irq <= Std_Logic_Vector'(A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(epcs_flash_controller_0_epcs_control_port_irq_from_sa) & A_ToStdLogicVector(clk90Meg_jtag_uart_0_avalon_jtag_slave_irq_from_sa) & A_ToStdLogicVector(clk90Meg_system_timer_s1_irq_from_sa) & A_ToStdLogicVector(clk90Meg_OpenMAC_0_REG_irq_from_sa) & A_ToStdLogicVector(clk90Meg_OpenMAC_0_CMP_irq_from_sa));
  --OpenMAC_0_REG_irq_from_sa from clk50Meg to clk90Meg
  OpenMAC_0_REG_irq_from_sa_clock_crossing_pcp_cpu_data_master : OpenMAC_0_REG_irq_from_sa_clock_crossing_pcp_cpu_data_master_module
    port map(
      data_out => clk90Meg_OpenMAC_0_REG_irq_from_sa,
      clk => clk90Meg,
      data_in => OpenMAC_0_REG_irq_from_sa,
      reset_n => clk90Meg_reset_n
    );


  --optimize select-logic by passing only those address bits which matter.
  internal_pcp_cpu_data_master_address_to_slave <= Std_Logic_Vector'(pcp_cpu_data_master_address(25 DOWNTO 24) & A_ToStdLogicVector(std_logic'('0')) & pcp_cpu_data_master_address(22 DOWNTO 0));
  --pcp_cpu/data_master readdata mux, which is an e_mux
  pcp_cpu_data_master_readdata <= (((((((((((((A_REP(NOT pcp_cpu_data_master_requests_OpenMAC_0_iBuf, 32) OR OpenMAC_0_iBuf_readdata_from_sa)) AND ((A_REP(NOT pcp_cpu_data_master_requests_clock_crossing_0_s1, 32) OR registered_pcp_cpu_data_master_readdata))) AND ((A_REP(NOT pcp_cpu_data_master_requests_cnApi_Av2Av_0_pcp, 32) OR cnApi_Av2Av_0_pcp_readdata_from_sa))) AND ((A_REP(NOT pcp_cpu_data_master_requests_epcs_flash_controller_0_epcs_control_port, 32) OR epcs_flash_controller_0_epcs_control_port_readdata_from_sa))) AND ((A_REP(NOT pcp_cpu_data_master_requests_niosII_openMac_clock_0_in, 32) OR registered_pcp_cpu_data_master_readdata))) AND ((A_REP(NOT pcp_cpu_data_master_requests_niosII_openMac_clock_1_in, 32) OR registered_pcp_cpu_data_master_readdata))) AND ((A_REP(NOT pcp_cpu_data_master_requests_niosII_openMac_clock_2_in, 32) OR registered_pcp_cpu_data_master_readdata))) AND ((A_REP(NOT pcp_cpu_data_master_requests_niosII_openMac_clock_3_in, 32) OR registered_pcp_cpu_data_master_readdata))) AND ((A_REP(NOT pcp_cpu_data_master_requests_niosII_openMac_clock_4_in, 32) OR registered_pcp_cpu_data_master_readdata))) AND ((A_REP(NOT pcp_cpu_data_master_requests_onchip_memory_0_s1, 32) OR onchip_memory_0_s1_readdata_from_sa))) AND ((A_REP(NOT pcp_cpu_data_master_requests_pcp_cpu_jtag_debug_module, 32) OR pcp_cpu_jtag_debug_module_readdata_from_sa))) AND ((A_REP(NOT pcp_cpu_data_master_requests_DBC3C40_SRAM_0_avalon_tristate_slave, 32) OR Std_Logic_Vector'(incoming_tri_state_bridge_0_data(15 DOWNTO 0) & dbs_16_reg_segment_0)))) AND ((A_REP(NOT pcp_cpu_data_master_requests_cfi_flash_0_s1, 32) OR Std_Logic_Vector'(incoming_tri_state_bridge_0_data_with_Xs_converted_to_0(15 DOWNTO 0) & dbs_16_reg_segment_0)));
  --actual waitrequest port, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      internal_pcp_cpu_data_master_waitrequest <= Vector_To_Std_Logic(NOT std_logic_vector'("00000000000000000000000000000000"));
    elsif clk'event and clk = '1' then
      internal_pcp_cpu_data_master_waitrequest <= Vector_To_Std_Logic(NOT (A_WE_StdLogicVector((std_logic'((NOT ((pcp_cpu_data_master_read OR pcp_cpu_data_master_write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pcp_cpu_data_master_run AND internal_pcp_cpu_data_master_waitrequest))))))));
    end if;

  end process;

  --unpredictable registered wait state incoming data, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      registered_pcp_cpu_data_master_readdata <= std_logic_vector'("00000000000000000000000000000000");
    elsif clk'event and clk = '1' then
      registered_pcp_cpu_data_master_readdata <= p1_registered_pcp_cpu_data_master_readdata;
    end if;

  end process;

  --registered readdata mux, which is an e_mux
  p1_registered_pcp_cpu_data_master_readdata <= ((((((A_REP(NOT pcp_cpu_data_master_requests_clock_crossing_0_s1, 32) OR clock_crossing_0_s1_readdata_from_sa)) AND ((A_REP(NOT pcp_cpu_data_master_requests_niosII_openMac_clock_0_in, 32) OR niosII_openMac_clock_0_in_readdata_from_sa))) AND ((A_REP(NOT pcp_cpu_data_master_requests_niosII_openMac_clock_1_in, 32) OR niosII_openMac_clock_1_in_readdata_from_sa))) AND ((A_REP(NOT pcp_cpu_data_master_requests_niosII_openMac_clock_2_in, 32) OR Std_Logic_Vector'(niosII_openMac_clock_2_in_readdata_from_sa(15 DOWNTO 0) & dbs_16_reg_segment_0)))) AND ((A_REP(NOT pcp_cpu_data_master_requests_niosII_openMac_clock_3_in, 32) OR niosII_openMac_clock_3_in_readdata_from_sa))) AND ((A_REP(NOT pcp_cpu_data_master_requests_niosII_openMac_clock_4_in, 32) OR niosII_openMac_clock_4_in_readdata_from_sa));
  --jtag_uart_0_avalon_jtag_slave_irq_from_sa from clk50Meg to clk90Meg
  jtag_uart_0_avalon_jtag_slave_irq_from_sa_clock_crossing_pcp_cpu_data_master : jtag_uart_0_avalon_jtag_slave_irq_from_sa_clock_crossing_pcp_cpu_data_master_module
    port map(
      data_out => clk90Meg_jtag_uart_0_avalon_jtag_slave_irq_from_sa,
      clk => clk90Meg,
      data_in => jtag_uart_0_avalon_jtag_slave_irq_from_sa,
      reset_n => clk90Meg_reset_n
    );


  --no_byte_enables_and_last_term, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      internal_pcp_cpu_data_master_no_byte_enables_and_last_term <= std_logic'('0');
    elsif clk'event and clk = '1' then
      internal_pcp_cpu_data_master_no_byte_enables_and_last_term <= last_dbs_term_and_run;
    end if;

  end process;

  --compute the last dbs term, which is an e_mux
  last_dbs_term_and_run <= A_WE_StdLogic((std_logic'((pcp_cpu_data_master_requests_niosII_openMac_clock_2_in)) = '1'), (((to_std_logic(((internal_pcp_cpu_data_master_dbs_address = std_logic_vector'("10")))) AND pcp_cpu_data_master_write) AND NOT(or_reduce(pcp_cpu_data_master_byteenable_niosII_openMac_clock_2_in)))), A_WE_StdLogic((std_logic'((pcp_cpu_data_master_requests_DBC3C40_SRAM_0_avalon_tristate_slave)) = '1'), (((to_std_logic(((internal_pcp_cpu_data_master_dbs_address = std_logic_vector'("10")))) AND pcp_cpu_data_master_write) AND NOT(or_reduce(pcp_cpu_data_master_byteenable_DBC3C40_SRAM_0_avalon_tristate_slave)))), (((to_std_logic(((internal_pcp_cpu_data_master_dbs_address = std_logic_vector'("10")))) AND pcp_cpu_data_master_write) AND NOT(or_reduce(pcp_cpu_data_master_byteenable_cfi_flash_0_s1))))));
  --pre dbs count enable, which is an e_mux
  pre_dbs_count_enable <= Vector_To_Std_Logic((((((((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((((NOT internal_pcp_cpu_data_master_no_byte_enables_and_last_term) AND pcp_cpu_data_master_requests_niosII_openMac_clock_2_in) AND pcp_cpu_data_master_write) AND NOT(or_reduce(pcp_cpu_data_master_byteenable_niosII_openMac_clock_2_in))))))) OR (((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((pcp_cpu_data_master_granted_niosII_openMac_clock_2_in AND pcp_cpu_data_master_read)))) AND std_logic_vector'("00000000000000000000000000000001")) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT niosII_openMac_clock_2_in_waitrequest_from_sa)))))) OR (((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((pcp_cpu_data_master_granted_niosII_openMac_clock_2_in AND pcp_cpu_data_master_write)))) AND std_logic_vector'("00000000000000000000000000000001")) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT niosII_openMac_clock_2_in_waitrequest_from_sa)))))) OR (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((((NOT internal_pcp_cpu_data_master_no_byte_enables_and_last_term) AND pcp_cpu_data_master_requests_DBC3C40_SRAM_0_avalon_tristate_slave) AND pcp_cpu_data_master_write) AND NOT(or_reduce(pcp_cpu_data_master_byteenable_DBC3C40_SRAM_0_avalon_tristate_slave)))))))) OR (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((((NOT internal_pcp_cpu_data_master_no_byte_enables_and_last_term) AND pcp_cpu_data_master_requests_cfi_flash_0_s1) AND pcp_cpu_data_master_write) AND NOT(or_reduce(pcp_cpu_data_master_byteenable_cfi_flash_0_s1)))))))) OR (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pcp_cpu_data_master_read_data_valid_DBC3C40_SRAM_0_avalon_tristate_slave)))) OR (((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((pcp_cpu_data_master_granted_DBC3C40_SRAM_0_avalon_tristate_slave AND pcp_cpu_data_master_write)))) AND std_logic_vector'("00000000000000000000000000000001")) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((DBC3C40_SRAM_0_avalon_tristate_slave_wait_counter_eq_0 AND NOT d1_tri_state_bridge_0_avalon_slave_end_xfer)))))))) OR (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pcp_cpu_data_master_read_data_valid_cfi_flash_0_s1)))) OR (((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((pcp_cpu_data_master_granted_cfi_flash_0_s1 AND pcp_cpu_data_master_write)))) AND std_logic_vector'("00000000000000000000000000000001")) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cfi_flash_0_s1_wait_counter_eq_0 AND NOT d1_tri_state_bridge_0_avalon_slave_end_xfer)))))))));
  --input to dbs-16 stored 0, which is an e_mux
  p1_dbs_16_reg_segment_0 <= A_WE_StdLogicVector((std_logic'((pcp_cpu_data_master_requests_niosII_openMac_clock_2_in)) = '1'), niosII_openMac_clock_2_in_readdata_from_sa, A_WE_StdLogicVector((std_logic'((pcp_cpu_data_master_requests_DBC3C40_SRAM_0_avalon_tristate_slave)) = '1'), incoming_tri_state_bridge_0_data, incoming_tri_state_bridge_0_data_with_Xs_converted_to_0));
  --dbs register for dbs-16 segment 0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      dbs_16_reg_segment_0 <= std_logic_vector'("0000000000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((dbs_count_enable AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((internal_pcp_cpu_data_master_dbs_address(1))))) = std_logic_vector'("00000000000000000000000000000000")))))) = '1' then 
        dbs_16_reg_segment_0 <= p1_dbs_16_reg_segment_0;
      end if;
    end if;

  end process;

  --mux write dbs 1, which is an e_mux
  pcp_cpu_data_master_dbs_write_16 <= A_WE_StdLogicVector((std_logic'((internal_pcp_cpu_data_master_dbs_address(1))) = '1'), pcp_cpu_data_master_writedata(31 DOWNTO 16), A_WE_StdLogicVector((std_logic'((NOT (internal_pcp_cpu_data_master_dbs_address(1)))) = '1'), pcp_cpu_data_master_writedata(15 DOWNTO 0), A_WE_StdLogicVector((std_logic'((internal_pcp_cpu_data_master_dbs_address(1))) = '1'), pcp_cpu_data_master_writedata(31 DOWNTO 16), A_WE_StdLogicVector((std_logic'((NOT (internal_pcp_cpu_data_master_dbs_address(1)))) = '1'), pcp_cpu_data_master_writedata(15 DOWNTO 0), A_WE_StdLogicVector((std_logic'((internal_pcp_cpu_data_master_dbs_address(1))) = '1'), pcp_cpu_data_master_writedata(31 DOWNTO 16), pcp_cpu_data_master_writedata(15 DOWNTO 0))))));
  --dbs count increment, which is an e_mux
  pcp_cpu_data_master_dbs_increment <= A_EXT (A_WE_StdLogicVector((std_logic'((pcp_cpu_data_master_requests_niosII_openMac_clock_2_in)) = '1'), std_logic_vector'("00000000000000000000000000000010"), A_WE_StdLogicVector((std_logic'((pcp_cpu_data_master_requests_DBC3C40_SRAM_0_avalon_tristate_slave)) = '1'), std_logic_vector'("00000000000000000000000000000010"), A_WE_StdLogicVector((std_logic'((pcp_cpu_data_master_requests_cfi_flash_0_s1)) = '1'), std_logic_vector'("00000000000000000000000000000010"), std_logic_vector'("00000000000000000000000000000000")))), 2);
  --dbs counter overflow, which is an e_assign
  dbs_counter_overflow <= internal_pcp_cpu_data_master_dbs_address(1) AND NOT((next_dbs_address(1)));
  --next master address, which is an e_assign
  next_dbs_address <= A_EXT (((std_logic_vector'("0") & (internal_pcp_cpu_data_master_dbs_address)) + (std_logic_vector'("0") & (pcp_cpu_data_master_dbs_increment))), 2);
  --dbs count enable, which is an e_mux
  dbs_count_enable <= pre_dbs_count_enable AND (NOT ((pcp_cpu_data_master_requests_niosII_openMac_clock_2_in AND NOT internal_pcp_cpu_data_master_waitrequest)));
  --dbs counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      internal_pcp_cpu_data_master_dbs_address <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      if std_logic'(dbs_count_enable) = '1' then 
        internal_pcp_cpu_data_master_dbs_address <= next_dbs_address;
      end if;
    end if;

  end process;

  --system_timer_s1_irq_from_sa from clk50Meg to clk90Meg
  system_timer_s1_irq_from_sa_clock_crossing_pcp_cpu_data_master : system_timer_s1_irq_from_sa_clock_crossing_pcp_cpu_data_master_module
    port map(
      data_out => clk90Meg_system_timer_s1_irq_from_sa,
      clk => clk90Meg,
      data_in => system_timer_s1_irq_from_sa,
      reset_n => clk90Meg_reset_n
    );


  --vhdl renameroo for output signals
  pcp_cpu_data_master_address_to_slave <= internal_pcp_cpu_data_master_address_to_slave;
  --vhdl renameroo for output signals
  pcp_cpu_data_master_dbs_address <= internal_pcp_cpu_data_master_dbs_address;
  --vhdl renameroo for output signals
  pcp_cpu_data_master_no_byte_enables_and_last_term <= internal_pcp_cpu_data_master_no_byte_enables_and_last_term;
  --vhdl renameroo for output signals
  pcp_cpu_data_master_waitrequest <= internal_pcp_cpu_data_master_waitrequest;

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity pcp_cpu_instruction_master_arbitrator is 
        port (
              -- inputs:
                 signal DBC3C40_SRAM_0_avalon_tristate_slave_wait_counter_eq_0 : IN STD_LOGIC;
                 signal cfi_flash_0_s1_wait_counter_eq_0 : IN STD_LOGIC;
                 signal cfi_flash_0_s1_wait_counter_eq_1 : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal d1_epcs_flash_controller_0_epcs_control_port_end_xfer : IN STD_LOGIC;
                 signal d1_onchip_memory_0_s1_end_xfer : IN STD_LOGIC;
                 signal d1_pcp_cpu_jtag_debug_module_end_xfer : IN STD_LOGIC;
                 signal d1_tri_state_bridge_0_avalon_slave_end_xfer : IN STD_LOGIC;
                 signal epcs_flash_controller_0_epcs_control_port_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal incoming_tri_state_bridge_0_data : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal onchip_memory_0_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal pcp_cpu_instruction_master_address : IN STD_LOGIC_VECTOR (25 DOWNTO 0);
                 signal pcp_cpu_instruction_master_granted_DBC3C40_SRAM_0_avalon_tristate_slave : IN STD_LOGIC;
                 signal pcp_cpu_instruction_master_granted_cfi_flash_0_s1 : IN STD_LOGIC;
                 signal pcp_cpu_instruction_master_granted_epcs_flash_controller_0_epcs_control_port : IN STD_LOGIC;
                 signal pcp_cpu_instruction_master_granted_onchip_memory_0_s1 : IN STD_LOGIC;
                 signal pcp_cpu_instruction_master_granted_pcp_cpu_jtag_debug_module : IN STD_LOGIC;
                 signal pcp_cpu_instruction_master_qualified_request_DBC3C40_SRAM_0_avalon_tristate_slave : IN STD_LOGIC;
                 signal pcp_cpu_instruction_master_qualified_request_cfi_flash_0_s1 : IN STD_LOGIC;
                 signal pcp_cpu_instruction_master_qualified_request_epcs_flash_controller_0_epcs_control_port : IN STD_LOGIC;
                 signal pcp_cpu_instruction_master_qualified_request_onchip_memory_0_s1 : IN STD_LOGIC;
                 signal pcp_cpu_instruction_master_qualified_request_pcp_cpu_jtag_debug_module : IN STD_LOGIC;
                 signal pcp_cpu_instruction_master_read : IN STD_LOGIC;
                 signal pcp_cpu_instruction_master_read_data_valid_DBC3C40_SRAM_0_avalon_tristate_slave : IN STD_LOGIC;
                 signal pcp_cpu_instruction_master_read_data_valid_cfi_flash_0_s1 : IN STD_LOGIC;
                 signal pcp_cpu_instruction_master_read_data_valid_epcs_flash_controller_0_epcs_control_port : IN STD_LOGIC;
                 signal pcp_cpu_instruction_master_read_data_valid_onchip_memory_0_s1 : IN STD_LOGIC;
                 signal pcp_cpu_instruction_master_read_data_valid_pcp_cpu_jtag_debug_module : IN STD_LOGIC;
                 signal pcp_cpu_instruction_master_requests_DBC3C40_SRAM_0_avalon_tristate_slave : IN STD_LOGIC;
                 signal pcp_cpu_instruction_master_requests_cfi_flash_0_s1 : IN STD_LOGIC;
                 signal pcp_cpu_instruction_master_requests_epcs_flash_controller_0_epcs_control_port : IN STD_LOGIC;
                 signal pcp_cpu_instruction_master_requests_onchip_memory_0_s1 : IN STD_LOGIC;
                 signal pcp_cpu_instruction_master_requests_pcp_cpu_jtag_debug_module : IN STD_LOGIC;
                 signal pcp_cpu_jtag_debug_module_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal pcp_cpu_instruction_master_address_to_slave : OUT STD_LOGIC_VECTOR (25 DOWNTO 0);
                 signal pcp_cpu_instruction_master_dbs_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal pcp_cpu_instruction_master_latency_counter : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal pcp_cpu_instruction_master_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal pcp_cpu_instruction_master_readdatavalid : OUT STD_LOGIC;
                 signal pcp_cpu_instruction_master_waitrequest : OUT STD_LOGIC
              );
end entity pcp_cpu_instruction_master_arbitrator;


architecture europa of pcp_cpu_instruction_master_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal dbs_count_enable :  STD_LOGIC;
                signal dbs_counter_overflow :  STD_LOGIC;
                signal dbs_latent_16_reg_segment_0 :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal dbs_rdv_count_enable :  STD_LOGIC;
                signal dbs_rdv_counter_overflow :  STD_LOGIC;
                signal internal_pcp_cpu_instruction_master_address_to_slave :  STD_LOGIC_VECTOR (25 DOWNTO 0);
                signal internal_pcp_cpu_instruction_master_dbs_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal internal_pcp_cpu_instruction_master_latency_counter :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal internal_pcp_cpu_instruction_master_waitrequest :  STD_LOGIC;
                signal latency_load_value :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal next_dbs_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal p1_dbs_latent_16_reg_segment_0 :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal p1_pcp_cpu_instruction_master_latency_counter :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal pcp_cpu_instruction_master_address_last_time :  STD_LOGIC_VECTOR (25 DOWNTO 0);
                signal pcp_cpu_instruction_master_dbs_increment :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal pcp_cpu_instruction_master_dbs_rdv_counter :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal pcp_cpu_instruction_master_dbs_rdv_counter_inc :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal pcp_cpu_instruction_master_is_granted_some_slave :  STD_LOGIC;
                signal pcp_cpu_instruction_master_next_dbs_rdv_counter :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal pcp_cpu_instruction_master_read_but_no_slave_selected :  STD_LOGIC;
                signal pcp_cpu_instruction_master_read_last_time :  STD_LOGIC;
                signal pcp_cpu_instruction_master_run :  STD_LOGIC;
                signal pre_dbs_count_enable :  STD_LOGIC;
                signal pre_flush_pcp_cpu_instruction_master_readdatavalid :  STD_LOGIC;
                signal r_0 :  STD_LOGIC;
                signal r_1 :  STD_LOGIC;
                signal r_2 :  STD_LOGIC;

begin

  --r_0 master_run cascaded wait assignment, which is an e_assign
  r_0 <= Vector_To_Std_Logic((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pcp_cpu_instruction_master_qualified_request_epcs_flash_controller_0_epcs_control_port OR NOT pcp_cpu_instruction_master_requests_epcs_flash_controller_0_epcs_control_port)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pcp_cpu_instruction_master_granted_epcs_flash_controller_0_epcs_control_port OR NOT pcp_cpu_instruction_master_qualified_request_epcs_flash_controller_0_epcs_control_port)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT pcp_cpu_instruction_master_qualified_request_epcs_flash_controller_0_epcs_control_port OR NOT (pcp_cpu_instruction_master_read))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT d1_epcs_flash_controller_0_epcs_control_port_end_xfer)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((pcp_cpu_instruction_master_read))))))))));
  --cascaded wait assignment, which is an e_assign
  pcp_cpu_instruction_master_run <= (r_0 AND r_1) AND r_2;
  --r_1 master_run cascaded wait assignment, which is an e_assign
  r_1 <= Vector_To_Std_Logic((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pcp_cpu_instruction_master_qualified_request_onchip_memory_0_s1 OR NOT pcp_cpu_instruction_master_requests_onchip_memory_0_s1)))))));
  --r_2 master_run cascaded wait assignment, which is an e_assign
  r_2 <= Vector_To_Std_Logic((((((((((((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pcp_cpu_instruction_master_granted_onchip_memory_0_s1 OR NOT pcp_cpu_instruction_master_qualified_request_onchip_memory_0_s1))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT pcp_cpu_instruction_master_qualified_request_onchip_memory_0_s1 OR NOT pcp_cpu_instruction_master_read)))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pcp_cpu_instruction_master_read)))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pcp_cpu_instruction_master_qualified_request_pcp_cpu_jtag_debug_module OR NOT pcp_cpu_instruction_master_requests_pcp_cpu_jtag_debug_module)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pcp_cpu_instruction_master_granted_pcp_cpu_jtag_debug_module OR NOT pcp_cpu_instruction_master_qualified_request_pcp_cpu_jtag_debug_module)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT pcp_cpu_instruction_master_qualified_request_pcp_cpu_jtag_debug_module OR NOT pcp_cpu_instruction_master_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT d1_pcp_cpu_jtag_debug_module_end_xfer)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pcp_cpu_instruction_master_read)))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pcp_cpu_instruction_master_qualified_request_DBC3C40_SRAM_0_avalon_tristate_slave OR NOT pcp_cpu_instruction_master_requests_DBC3C40_SRAM_0_avalon_tristate_slave)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pcp_cpu_instruction_master_qualified_request_cfi_flash_0_s1 OR NOT pcp_cpu_instruction_master_requests_cfi_flash_0_s1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pcp_cpu_instruction_master_granted_DBC3C40_SRAM_0_avalon_tristate_slave OR NOT pcp_cpu_instruction_master_qualified_request_DBC3C40_SRAM_0_avalon_tristate_slave)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pcp_cpu_instruction_master_granted_cfi_flash_0_s1 OR NOT pcp_cpu_instruction_master_qualified_request_cfi_flash_0_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT pcp_cpu_instruction_master_qualified_request_DBC3C40_SRAM_0_avalon_tristate_slave OR NOT pcp_cpu_instruction_master_read)))) OR ((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((DBC3C40_SRAM_0_avalon_tristate_slave_wait_counter_eq_0 AND NOT d1_tri_state_bridge_0_avalon_slave_end_xfer)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((internal_pcp_cpu_instruction_master_dbs_address(1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pcp_cpu_instruction_master_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT pcp_cpu_instruction_master_qualified_request_cfi_flash_0_s1 OR NOT pcp_cpu_instruction_master_read)))) OR ((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cfi_flash_0_s1_wait_counter_eq_0 AND NOT d1_tri_state_bridge_0_avalon_slave_end_xfer)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((internal_pcp_cpu_instruction_master_dbs_address(1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pcp_cpu_instruction_master_read)))))))));
  --optimize select-logic by passing only those address bits which matter.
  internal_pcp_cpu_instruction_master_address_to_slave <= Std_Logic_Vector'(A_ToStdLogicVector(pcp_cpu_instruction_master_address(25)) & std_logic_vector'("00") & pcp_cpu_instruction_master_address(22 DOWNTO 0));
  --pcp_cpu_instruction_master_read_but_no_slave_selected assignment, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pcp_cpu_instruction_master_read_but_no_slave_selected <= std_logic'('0');
    elsif clk'event and clk = '1' then
      pcp_cpu_instruction_master_read_but_no_slave_selected <= (pcp_cpu_instruction_master_read AND pcp_cpu_instruction_master_run) AND NOT pcp_cpu_instruction_master_is_granted_some_slave;
    end if;

  end process;

  --some slave is getting selected, which is an e_mux
  pcp_cpu_instruction_master_is_granted_some_slave <= (((pcp_cpu_instruction_master_granted_epcs_flash_controller_0_epcs_control_port OR pcp_cpu_instruction_master_granted_onchip_memory_0_s1) OR pcp_cpu_instruction_master_granted_pcp_cpu_jtag_debug_module) OR pcp_cpu_instruction_master_granted_DBC3C40_SRAM_0_avalon_tristate_slave) OR pcp_cpu_instruction_master_granted_cfi_flash_0_s1;
  --latent slave read data valids which may be flushed, which is an e_mux
  pre_flush_pcp_cpu_instruction_master_readdatavalid <= (pcp_cpu_instruction_master_read_data_valid_onchip_memory_0_s1 OR ((pcp_cpu_instruction_master_read_data_valid_DBC3C40_SRAM_0_avalon_tristate_slave AND dbs_rdv_counter_overflow))) OR ((pcp_cpu_instruction_master_read_data_valid_cfi_flash_0_s1 AND dbs_rdv_counter_overflow));
  --latent slave read data valid which is not flushed, which is an e_mux
  pcp_cpu_instruction_master_readdatavalid <= ((((((((((pcp_cpu_instruction_master_read_but_no_slave_selected OR pre_flush_pcp_cpu_instruction_master_readdatavalid) OR pcp_cpu_instruction_master_read_data_valid_epcs_flash_controller_0_epcs_control_port) OR pcp_cpu_instruction_master_read_but_no_slave_selected) OR pre_flush_pcp_cpu_instruction_master_readdatavalid) OR pcp_cpu_instruction_master_read_but_no_slave_selected) OR pre_flush_pcp_cpu_instruction_master_readdatavalid) OR pcp_cpu_instruction_master_read_data_valid_pcp_cpu_jtag_debug_module) OR pcp_cpu_instruction_master_read_but_no_slave_selected) OR pre_flush_pcp_cpu_instruction_master_readdatavalid) OR pcp_cpu_instruction_master_read_but_no_slave_selected) OR pre_flush_pcp_cpu_instruction_master_readdatavalid;
  --pcp_cpu/instruction_master readdata mux, which is an e_mux
  pcp_cpu_instruction_master_readdata <= (((((A_REP(NOT ((pcp_cpu_instruction_master_qualified_request_epcs_flash_controller_0_epcs_control_port AND pcp_cpu_instruction_master_read)) , 32) OR epcs_flash_controller_0_epcs_control_port_readdata_from_sa)) AND ((A_REP(NOT pcp_cpu_instruction_master_read_data_valid_onchip_memory_0_s1, 32) OR onchip_memory_0_s1_readdata_from_sa))) AND ((A_REP(NOT ((pcp_cpu_instruction_master_qualified_request_pcp_cpu_jtag_debug_module AND pcp_cpu_instruction_master_read)) , 32) OR pcp_cpu_jtag_debug_module_readdata_from_sa))) AND ((A_REP(NOT pcp_cpu_instruction_master_read_data_valid_DBC3C40_SRAM_0_avalon_tristate_slave, 32) OR Std_Logic_Vector'(incoming_tri_state_bridge_0_data(15 DOWNTO 0) & dbs_latent_16_reg_segment_0)))) AND ((A_REP(NOT pcp_cpu_instruction_master_read_data_valid_cfi_flash_0_s1, 32) OR Std_Logic_Vector'(incoming_tri_state_bridge_0_data(15 DOWNTO 0) & dbs_latent_16_reg_segment_0)));
  --actual waitrequest port, which is an e_assign
  internal_pcp_cpu_instruction_master_waitrequest <= NOT pcp_cpu_instruction_master_run;
  --latent max counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      internal_pcp_cpu_instruction_master_latency_counter <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      internal_pcp_cpu_instruction_master_latency_counter <= p1_pcp_cpu_instruction_master_latency_counter;
    end if;

  end process;

  --latency counter load mux, which is an e_mux
  p1_pcp_cpu_instruction_master_latency_counter <= A_EXT (A_WE_StdLogicVector((std_logic'(((pcp_cpu_instruction_master_run AND pcp_cpu_instruction_master_read))) = '1'), (std_logic_vector'("0000000000000000000000000000000") & (latency_load_value)), A_WE_StdLogicVector((((internal_pcp_cpu_instruction_master_latency_counter)) /= std_logic_vector'("00")), ((std_logic_vector'("0000000000000000000000000000000") & (internal_pcp_cpu_instruction_master_latency_counter)) - std_logic_vector'("000000000000000000000000000000001")), std_logic_vector'("000000000000000000000000000000000"))), 2);
  --read latency load values, which is an e_mux
  latency_load_value <= A_EXT ((((((std_logic_vector'("000000000000000000000000000000") & (A_REP(pcp_cpu_instruction_master_requests_onchip_memory_0_s1, 2))) AND std_logic_vector'("00000000000000000000000000000001"))) OR (((std_logic_vector'("000000000000000000000000000000") & (A_REP(pcp_cpu_instruction_master_requests_DBC3C40_SRAM_0_avalon_tristate_slave, 2))) AND std_logic_vector'("00000000000000000000000000000010")))) OR (((std_logic_vector'("000000000000000000000000000000") & (A_REP(pcp_cpu_instruction_master_requests_cfi_flash_0_s1, 2))) AND std_logic_vector'("00000000000000000000000000000010")))), 2);
  --input to latent dbs-16 stored 0, which is an e_mux
  p1_dbs_latent_16_reg_segment_0 <= A_WE_StdLogicVector((std_logic'((pcp_cpu_instruction_master_read_data_valid_DBC3C40_SRAM_0_avalon_tristate_slave)) = '1'), incoming_tri_state_bridge_0_data, incoming_tri_state_bridge_0_data);
  --dbs register for latent dbs-16 segment 0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      dbs_latent_16_reg_segment_0 <= std_logic_vector'("0000000000000000");
    elsif clk'event and clk = '1' then
      if std_logic'((dbs_rdv_count_enable AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((pcp_cpu_instruction_master_dbs_rdv_counter(1))))) = std_logic_vector'("00000000000000000000000000000000")))))) = '1' then 
        dbs_latent_16_reg_segment_0 <= p1_dbs_latent_16_reg_segment_0;
      end if;
    end if;

  end process;

  --dbs count increment, which is an e_mux
  pcp_cpu_instruction_master_dbs_increment <= A_EXT (A_WE_StdLogicVector((std_logic'((pcp_cpu_instruction_master_requests_DBC3C40_SRAM_0_avalon_tristate_slave)) = '1'), std_logic_vector'("00000000000000000000000000000010"), A_WE_StdLogicVector((std_logic'((pcp_cpu_instruction_master_requests_cfi_flash_0_s1)) = '1'), std_logic_vector'("00000000000000000000000000000010"), std_logic_vector'("00000000000000000000000000000000"))), 2);
  --dbs counter overflow, which is an e_assign
  dbs_counter_overflow <= internal_pcp_cpu_instruction_master_dbs_address(1) AND NOT((next_dbs_address(1)));
  --next master address, which is an e_assign
  next_dbs_address <= A_EXT (((std_logic_vector'("0") & (internal_pcp_cpu_instruction_master_dbs_address)) + (std_logic_vector'("0") & (pcp_cpu_instruction_master_dbs_increment))), 2);
  --dbs count enable, which is an e_mux
  dbs_count_enable <= pre_dbs_count_enable;
  --dbs counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      internal_pcp_cpu_instruction_master_dbs_address <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      if std_logic'(dbs_count_enable) = '1' then 
        internal_pcp_cpu_instruction_master_dbs_address <= next_dbs_address;
      end if;
    end if;

  end process;

  --p1 dbs rdv counter, which is an e_assign
  pcp_cpu_instruction_master_next_dbs_rdv_counter <= A_EXT (((std_logic_vector'("0") & (pcp_cpu_instruction_master_dbs_rdv_counter)) + (std_logic_vector'("0") & (pcp_cpu_instruction_master_dbs_rdv_counter_inc))), 2);
  --pcp_cpu_instruction_master_rdv_inc_mux, which is an e_mux
  pcp_cpu_instruction_master_dbs_rdv_counter_inc <= A_EXT (A_WE_StdLogicVector((std_logic'((pcp_cpu_instruction_master_read_data_valid_DBC3C40_SRAM_0_avalon_tristate_slave)) = '1'), std_logic_vector'("00000000000000000000000000000010"), std_logic_vector'("00000000000000000000000000000010")), 2);
  --master any slave rdv, which is an e_mux
  dbs_rdv_count_enable <= pcp_cpu_instruction_master_read_data_valid_DBC3C40_SRAM_0_avalon_tristate_slave OR pcp_cpu_instruction_master_read_data_valid_cfi_flash_0_s1;
  --dbs rdv counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pcp_cpu_instruction_master_dbs_rdv_counter <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      if std_logic'(dbs_rdv_count_enable) = '1' then 
        pcp_cpu_instruction_master_dbs_rdv_counter <= pcp_cpu_instruction_master_next_dbs_rdv_counter;
      end if;
    end if;

  end process;

  --dbs rdv counter overflow, which is an e_assign
  dbs_rdv_counter_overflow <= pcp_cpu_instruction_master_dbs_rdv_counter(1) AND NOT pcp_cpu_instruction_master_next_dbs_rdv_counter(1);
  --pre dbs count enable, which is an e_mux
  pre_dbs_count_enable <= Vector_To_Std_Logic(((((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((pcp_cpu_instruction_master_granted_DBC3C40_SRAM_0_avalon_tristate_slave AND pcp_cpu_instruction_master_read)))) AND std_logic_vector'("00000000000000000000000000000001")) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((DBC3C40_SRAM_0_avalon_tristate_slave_wait_counter_eq_0 AND NOT d1_tri_state_bridge_0_avalon_slave_end_xfer))))))) OR (((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((pcp_cpu_instruction_master_granted_cfi_flash_0_s1 AND pcp_cpu_instruction_master_read)))) AND std_logic_vector'("00000000000000000000000000000001")) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cfi_flash_0_s1_wait_counter_eq_0 AND NOT d1_tri_state_bridge_0_avalon_slave_end_xfer)))))))));
  --vhdl renameroo for output signals
  pcp_cpu_instruction_master_address_to_slave <= internal_pcp_cpu_instruction_master_address_to_slave;
  --vhdl renameroo for output signals
  pcp_cpu_instruction_master_dbs_address <= internal_pcp_cpu_instruction_master_dbs_address;
  --vhdl renameroo for output signals
  pcp_cpu_instruction_master_latency_counter <= internal_pcp_cpu_instruction_master_latency_counter;
  --vhdl renameroo for output signals
  pcp_cpu_instruction_master_waitrequest <= internal_pcp_cpu_instruction_master_waitrequest;
--synthesis translate_off
    --pcp_cpu_instruction_master_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        pcp_cpu_instruction_master_address_last_time <= std_logic_vector'("00000000000000000000000000");
      elsif clk'event and clk = '1' then
        pcp_cpu_instruction_master_address_last_time <= pcp_cpu_instruction_master_address;
      end if;

    end process;

    --pcp_cpu/instruction_master waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_pcp_cpu_instruction_master_waitrequest AND (pcp_cpu_instruction_master_read);
      end if;

    end process;

    --pcp_cpu_instruction_master_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line45 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((pcp_cpu_instruction_master_address /= pcp_cpu_instruction_master_address_last_time))))) = '1' then 
          write(write_line45, now);
          write(write_line45, string'(": "));
          write(write_line45, string'("pcp_cpu_instruction_master_address did not heed wait!!!"));
          write(output, write_line45.all);
          deallocate (write_line45);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --pcp_cpu_instruction_master_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        pcp_cpu_instruction_master_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        pcp_cpu_instruction_master_read_last_time <= pcp_cpu_instruction_master_read;
      end if;

    end process;

    --pcp_cpu_instruction_master_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line46 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(pcp_cpu_instruction_master_read) /= std_logic'(pcp_cpu_instruction_master_read_last_time)))))) = '1' then 
          write(write_line46, now);
          write(write_line46, string'(": "));
          write(write_line46, string'("pcp_cpu_instruction_master_read did not heed wait!!!"));
          write(output, write_line46.all);
          deallocate (write_line46);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity portconf_pio_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal clock_crossing_1_m1_address_to_slave : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal clock_crossing_1_m1_latency_counter : IN STD_LOGIC;
                 signal clock_crossing_1_m1_nativeaddress : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
                 signal clock_crossing_1_m1_read : IN STD_LOGIC;
                 signal clock_crossing_1_m1_write : IN STD_LOGIC;
                 signal clock_crossing_1_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal portconf_pio_s1_readdata : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal clock_crossing_1_m1_granted_portconf_pio_s1 : OUT STD_LOGIC;
                 signal clock_crossing_1_m1_qualified_request_portconf_pio_s1 : OUT STD_LOGIC;
                 signal clock_crossing_1_m1_read_data_valid_portconf_pio_s1 : OUT STD_LOGIC;
                 signal clock_crossing_1_m1_requests_portconf_pio_s1 : OUT STD_LOGIC;
                 signal d1_portconf_pio_s1_end_xfer : OUT STD_LOGIC;
                 signal portconf_pio_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal portconf_pio_s1_chipselect : OUT STD_LOGIC;
                 signal portconf_pio_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal portconf_pio_s1_reset_n : OUT STD_LOGIC;
                 signal portconf_pio_s1_write_n : OUT STD_LOGIC;
                 signal portconf_pio_s1_writedata : OUT STD_LOGIC_VECTOR (3 DOWNTO 0)
              );
end entity portconf_pio_s1_arbitrator;


architecture europa of portconf_pio_s1_arbitrator is
                signal clock_crossing_1_m1_arbiterlock :  STD_LOGIC;
                signal clock_crossing_1_m1_arbiterlock2 :  STD_LOGIC;
                signal clock_crossing_1_m1_continuerequest :  STD_LOGIC;
                signal clock_crossing_1_m1_saved_grant_portconf_pio_s1 :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_portconf_pio_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_clock_crossing_1_m1_granted_portconf_pio_s1 :  STD_LOGIC;
                signal internal_clock_crossing_1_m1_qualified_request_portconf_pio_s1 :  STD_LOGIC;
                signal internal_clock_crossing_1_m1_requests_portconf_pio_s1 :  STD_LOGIC;
                signal portconf_pio_s1_allgrants :  STD_LOGIC;
                signal portconf_pio_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal portconf_pio_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal portconf_pio_s1_any_continuerequest :  STD_LOGIC;
                signal portconf_pio_s1_arb_counter_enable :  STD_LOGIC;
                signal portconf_pio_s1_arb_share_counter :  STD_LOGIC;
                signal portconf_pio_s1_arb_share_counter_next_value :  STD_LOGIC;
                signal portconf_pio_s1_arb_share_set_values :  STD_LOGIC;
                signal portconf_pio_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal portconf_pio_s1_begins_xfer :  STD_LOGIC;
                signal portconf_pio_s1_end_xfer :  STD_LOGIC;
                signal portconf_pio_s1_firsttransfer :  STD_LOGIC;
                signal portconf_pio_s1_grant_vector :  STD_LOGIC;
                signal portconf_pio_s1_in_a_read_cycle :  STD_LOGIC;
                signal portconf_pio_s1_in_a_write_cycle :  STD_LOGIC;
                signal portconf_pio_s1_master_qreq_vector :  STD_LOGIC;
                signal portconf_pio_s1_non_bursting_master_requests :  STD_LOGIC;
                signal portconf_pio_s1_reg_firsttransfer :  STD_LOGIC;
                signal portconf_pio_s1_slavearbiterlockenable :  STD_LOGIC;
                signal portconf_pio_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal portconf_pio_s1_unreg_firsttransfer :  STD_LOGIC;
                signal portconf_pio_s1_waits_for_read :  STD_LOGIC;
                signal portconf_pio_s1_waits_for_write :  STD_LOGIC;
                signal wait_for_portconf_pio_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT portconf_pio_s1_end_xfer;
    end if;

  end process;

  portconf_pio_s1_begins_xfer <= NOT d1_reasons_to_wait AND (internal_clock_crossing_1_m1_qualified_request_portconf_pio_s1);
  --assign portconf_pio_s1_readdata_from_sa = portconf_pio_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  portconf_pio_s1_readdata_from_sa <= portconf_pio_s1_readdata;
  internal_clock_crossing_1_m1_requests_portconf_pio_s1 <= to_std_logic(((Std_Logic_Vector'(clock_crossing_1_m1_address_to_slave(7 DOWNTO 4) & std_logic_vector'("0000")) = std_logic_vector'("01110000")))) AND ((clock_crossing_1_m1_read OR clock_crossing_1_m1_write));
  --portconf_pio_s1_arb_share_counter set values, which is an e_mux
  portconf_pio_s1_arb_share_set_values <= std_logic'('1');
  --portconf_pio_s1_non_bursting_master_requests mux, which is an e_mux
  portconf_pio_s1_non_bursting_master_requests <= internal_clock_crossing_1_m1_requests_portconf_pio_s1;
  --portconf_pio_s1_any_bursting_master_saved_grant mux, which is an e_mux
  portconf_pio_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --portconf_pio_s1_arb_share_counter_next_value assignment, which is an e_assign
  portconf_pio_s1_arb_share_counter_next_value <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(portconf_pio_s1_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(portconf_pio_s1_arb_share_set_values))) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(portconf_pio_s1_arb_share_counter) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(portconf_pio_s1_arb_share_counter))) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))));
  --portconf_pio_s1_allgrants all slave grants, which is an e_mux
  portconf_pio_s1_allgrants <= portconf_pio_s1_grant_vector;
  --portconf_pio_s1_end_xfer assignment, which is an e_assign
  portconf_pio_s1_end_xfer <= NOT ((portconf_pio_s1_waits_for_read OR portconf_pio_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_portconf_pio_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_portconf_pio_s1 <= portconf_pio_s1_end_xfer AND (((NOT portconf_pio_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --portconf_pio_s1_arb_share_counter arbitration counter enable, which is an e_assign
  portconf_pio_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_portconf_pio_s1 AND portconf_pio_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_portconf_pio_s1 AND NOT portconf_pio_s1_non_bursting_master_requests));
  --portconf_pio_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      portconf_pio_s1_arb_share_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(portconf_pio_s1_arb_counter_enable) = '1' then 
        portconf_pio_s1_arb_share_counter <= portconf_pio_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --portconf_pio_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      portconf_pio_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((portconf_pio_s1_master_qreq_vector AND end_xfer_arb_share_counter_term_portconf_pio_s1)) OR ((end_xfer_arb_share_counter_term_portconf_pio_s1 AND NOT portconf_pio_s1_non_bursting_master_requests)))) = '1' then 
        portconf_pio_s1_slavearbiterlockenable <= portconf_pio_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --clock_crossing_1/m1 portconf_pio/s1 arbiterlock, which is an e_assign
  clock_crossing_1_m1_arbiterlock <= portconf_pio_s1_slavearbiterlockenable AND clock_crossing_1_m1_continuerequest;
  --portconf_pio_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  portconf_pio_s1_slavearbiterlockenable2 <= portconf_pio_s1_arb_share_counter_next_value;
  --clock_crossing_1/m1 portconf_pio/s1 arbiterlock2, which is an e_assign
  clock_crossing_1_m1_arbiterlock2 <= portconf_pio_s1_slavearbiterlockenable2 AND clock_crossing_1_m1_continuerequest;
  --portconf_pio_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  portconf_pio_s1_any_continuerequest <= std_logic'('1');
  --clock_crossing_1_m1_continuerequest continued request, which is an e_assign
  clock_crossing_1_m1_continuerequest <= std_logic'('1');
  internal_clock_crossing_1_m1_qualified_request_portconf_pio_s1 <= internal_clock_crossing_1_m1_requests_portconf_pio_s1 AND NOT ((clock_crossing_1_m1_read AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(clock_crossing_1_m1_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))))));
  --local readdatavalid clock_crossing_1_m1_read_data_valid_portconf_pio_s1, which is an e_mux
  clock_crossing_1_m1_read_data_valid_portconf_pio_s1 <= (internal_clock_crossing_1_m1_granted_portconf_pio_s1 AND clock_crossing_1_m1_read) AND NOT portconf_pio_s1_waits_for_read;
  --portconf_pio_s1_writedata mux, which is an e_mux
  portconf_pio_s1_writedata <= clock_crossing_1_m1_writedata (3 DOWNTO 0);
  --master is always granted when requested
  internal_clock_crossing_1_m1_granted_portconf_pio_s1 <= internal_clock_crossing_1_m1_qualified_request_portconf_pio_s1;
  --clock_crossing_1/m1 saved-grant portconf_pio/s1, which is an e_assign
  clock_crossing_1_m1_saved_grant_portconf_pio_s1 <= internal_clock_crossing_1_m1_requests_portconf_pio_s1;
  --allow new arb cycle for portconf_pio/s1, which is an e_assign
  portconf_pio_s1_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  portconf_pio_s1_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  portconf_pio_s1_master_qreq_vector <= std_logic'('1');
  --portconf_pio_s1_reset_n assignment, which is an e_assign
  portconf_pio_s1_reset_n <= reset_n;
  portconf_pio_s1_chipselect <= internal_clock_crossing_1_m1_granted_portconf_pio_s1;
  --portconf_pio_s1_firsttransfer first transaction, which is an e_assign
  portconf_pio_s1_firsttransfer <= A_WE_StdLogic((std_logic'(portconf_pio_s1_begins_xfer) = '1'), portconf_pio_s1_unreg_firsttransfer, portconf_pio_s1_reg_firsttransfer);
  --portconf_pio_s1_unreg_firsttransfer first transaction, which is an e_assign
  portconf_pio_s1_unreg_firsttransfer <= NOT ((portconf_pio_s1_slavearbiterlockenable AND portconf_pio_s1_any_continuerequest));
  --portconf_pio_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      portconf_pio_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(portconf_pio_s1_begins_xfer) = '1' then 
        portconf_pio_s1_reg_firsttransfer <= portconf_pio_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --portconf_pio_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  portconf_pio_s1_beginbursttransfer_internal <= portconf_pio_s1_begins_xfer;
  --~portconf_pio_s1_write_n assignment, which is an e_mux
  portconf_pio_s1_write_n <= NOT ((internal_clock_crossing_1_m1_granted_portconf_pio_s1 AND clock_crossing_1_m1_write));
  --portconf_pio_s1_address mux, which is an e_mux
  portconf_pio_s1_address <= clock_crossing_1_m1_nativeaddress (1 DOWNTO 0);
  --d1_portconf_pio_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_portconf_pio_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_portconf_pio_s1_end_xfer <= portconf_pio_s1_end_xfer;
    end if;

  end process;

  --portconf_pio_s1_waits_for_read in a cycle, which is an e_mux
  portconf_pio_s1_waits_for_read <= portconf_pio_s1_in_a_read_cycle AND portconf_pio_s1_begins_xfer;
  --portconf_pio_s1_in_a_read_cycle assignment, which is an e_assign
  portconf_pio_s1_in_a_read_cycle <= internal_clock_crossing_1_m1_granted_portconf_pio_s1 AND clock_crossing_1_m1_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= portconf_pio_s1_in_a_read_cycle;
  --portconf_pio_s1_waits_for_write in a cycle, which is an e_mux
  portconf_pio_s1_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(portconf_pio_s1_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --portconf_pio_s1_in_a_write_cycle assignment, which is an e_assign
  portconf_pio_s1_in_a_write_cycle <= internal_clock_crossing_1_m1_granted_portconf_pio_s1 AND clock_crossing_1_m1_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= portconf_pio_s1_in_a_write_cycle;
  wait_for_portconf_pio_s1_counter <= std_logic'('0');
  --vhdl renameroo for output signals
  clock_crossing_1_m1_granted_portconf_pio_s1 <= internal_clock_crossing_1_m1_granted_portconf_pio_s1;
  --vhdl renameroo for output signals
  clock_crossing_1_m1_qualified_request_portconf_pio_s1 <= internal_clock_crossing_1_m1_qualified_request_portconf_pio_s1;
  --vhdl renameroo for output signals
  clock_crossing_1_m1_requests_portconf_pio_s1 <= internal_clock_crossing_1_m1_requests_portconf_pio_s1;
--synthesis translate_off
    --portconf_pio/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity remote_update_cycloneiii_0_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal niosII_openMac_clock_4_out_address_to_slave : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal niosII_openMac_clock_4_out_nativeaddress : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
                 signal niosII_openMac_clock_4_out_read : IN STD_LOGIC;
                 signal niosII_openMac_clock_4_out_write : IN STD_LOGIC;
                 signal niosII_openMac_clock_4_out_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal remote_update_cycloneiii_0_s1_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal remote_update_cycloneiii_0_s1_waitrequest : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal d1_remote_update_cycloneiii_0_s1_end_xfer : OUT STD_LOGIC;
                 signal niosII_openMac_clock_4_out_granted_remote_update_cycloneiii_0_s1 : OUT STD_LOGIC;
                 signal niosII_openMac_clock_4_out_qualified_request_remote_update_cycloneiii_0_s1 : OUT STD_LOGIC;
                 signal niosII_openMac_clock_4_out_read_data_valid_remote_update_cycloneiii_0_s1 : OUT STD_LOGIC;
                 signal niosII_openMac_clock_4_out_requests_remote_update_cycloneiii_0_s1 : OUT STD_LOGIC;
                 signal remote_update_cycloneiii_0_s1_address : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
                 signal remote_update_cycloneiii_0_s1_chipselect : OUT STD_LOGIC;
                 signal remote_update_cycloneiii_0_s1_read : OUT STD_LOGIC;
                 signal remote_update_cycloneiii_0_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal remote_update_cycloneiii_0_s1_reset : OUT STD_LOGIC;
                 signal remote_update_cycloneiii_0_s1_waitrequest_from_sa : OUT STD_LOGIC;
                 signal remote_update_cycloneiii_0_s1_write : OUT STD_LOGIC;
                 signal remote_update_cycloneiii_0_s1_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
              );
end entity remote_update_cycloneiii_0_s1_arbitrator;


architecture europa of remote_update_cycloneiii_0_s1_arbitrator is
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_remote_update_cycloneiii_0_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_niosII_openMac_clock_4_out_granted_remote_update_cycloneiii_0_s1 :  STD_LOGIC;
                signal internal_niosII_openMac_clock_4_out_qualified_request_remote_update_cycloneiii_0_s1 :  STD_LOGIC;
                signal internal_niosII_openMac_clock_4_out_requests_remote_update_cycloneiii_0_s1 :  STD_LOGIC;
                signal internal_remote_update_cycloneiii_0_s1_waitrequest_from_sa :  STD_LOGIC;
                signal niosII_openMac_clock_4_out_arbiterlock :  STD_LOGIC;
                signal niosII_openMac_clock_4_out_arbiterlock2 :  STD_LOGIC;
                signal niosII_openMac_clock_4_out_continuerequest :  STD_LOGIC;
                signal niosII_openMac_clock_4_out_read_data_valid_remote_update_cycloneiii_0_s1_shift_register :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal niosII_openMac_clock_4_out_read_data_valid_remote_update_cycloneiii_0_s1_shift_register_in :  STD_LOGIC;
                signal niosII_openMac_clock_4_out_saved_grant_remote_update_cycloneiii_0_s1 :  STD_LOGIC;
                signal p1_niosII_openMac_clock_4_out_read_data_valid_remote_update_cycloneiii_0_s1_shift_register :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal remote_update_cycloneiii_0_s1_allgrants :  STD_LOGIC;
                signal remote_update_cycloneiii_0_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal remote_update_cycloneiii_0_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal remote_update_cycloneiii_0_s1_any_continuerequest :  STD_LOGIC;
                signal remote_update_cycloneiii_0_s1_arb_counter_enable :  STD_LOGIC;
                signal remote_update_cycloneiii_0_s1_arb_share_counter :  STD_LOGIC;
                signal remote_update_cycloneiii_0_s1_arb_share_counter_next_value :  STD_LOGIC;
                signal remote_update_cycloneiii_0_s1_arb_share_set_values :  STD_LOGIC;
                signal remote_update_cycloneiii_0_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal remote_update_cycloneiii_0_s1_begins_xfer :  STD_LOGIC;
                signal remote_update_cycloneiii_0_s1_end_xfer :  STD_LOGIC;
                signal remote_update_cycloneiii_0_s1_firsttransfer :  STD_LOGIC;
                signal remote_update_cycloneiii_0_s1_grant_vector :  STD_LOGIC;
                signal remote_update_cycloneiii_0_s1_in_a_read_cycle :  STD_LOGIC;
                signal remote_update_cycloneiii_0_s1_in_a_write_cycle :  STD_LOGIC;
                signal remote_update_cycloneiii_0_s1_master_qreq_vector :  STD_LOGIC;
                signal remote_update_cycloneiii_0_s1_non_bursting_master_requests :  STD_LOGIC;
                signal remote_update_cycloneiii_0_s1_reg_firsttransfer :  STD_LOGIC;
                signal remote_update_cycloneiii_0_s1_slavearbiterlockenable :  STD_LOGIC;
                signal remote_update_cycloneiii_0_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal remote_update_cycloneiii_0_s1_unreg_firsttransfer :  STD_LOGIC;
                signal remote_update_cycloneiii_0_s1_waits_for_read :  STD_LOGIC;
                signal remote_update_cycloneiii_0_s1_waits_for_write :  STD_LOGIC;
                signal wait_for_remote_update_cycloneiii_0_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT remote_update_cycloneiii_0_s1_end_xfer;
    end if;

  end process;

  remote_update_cycloneiii_0_s1_begins_xfer <= NOT d1_reasons_to_wait AND (internal_niosII_openMac_clock_4_out_qualified_request_remote_update_cycloneiii_0_s1);
  --assign remote_update_cycloneiii_0_s1_readdata_from_sa = remote_update_cycloneiii_0_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  remote_update_cycloneiii_0_s1_readdata_from_sa <= remote_update_cycloneiii_0_s1_readdata;
  internal_niosII_openMac_clock_4_out_requests_remote_update_cycloneiii_0_s1 <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((niosII_openMac_clock_4_out_read OR niosII_openMac_clock_4_out_write)))))));
  --assign remote_update_cycloneiii_0_s1_waitrequest_from_sa = remote_update_cycloneiii_0_s1_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_remote_update_cycloneiii_0_s1_waitrequest_from_sa <= remote_update_cycloneiii_0_s1_waitrequest;
  --remote_update_cycloneiii_0_s1_arb_share_counter set values, which is an e_mux
  remote_update_cycloneiii_0_s1_arb_share_set_values <= std_logic'('1');
  --remote_update_cycloneiii_0_s1_non_bursting_master_requests mux, which is an e_mux
  remote_update_cycloneiii_0_s1_non_bursting_master_requests <= internal_niosII_openMac_clock_4_out_requests_remote_update_cycloneiii_0_s1;
  --remote_update_cycloneiii_0_s1_any_bursting_master_saved_grant mux, which is an e_mux
  remote_update_cycloneiii_0_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --remote_update_cycloneiii_0_s1_arb_share_counter_next_value assignment, which is an e_assign
  remote_update_cycloneiii_0_s1_arb_share_counter_next_value <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(remote_update_cycloneiii_0_s1_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(remote_update_cycloneiii_0_s1_arb_share_set_values))) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(remote_update_cycloneiii_0_s1_arb_share_counter) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(remote_update_cycloneiii_0_s1_arb_share_counter))) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))));
  --remote_update_cycloneiii_0_s1_allgrants all slave grants, which is an e_mux
  remote_update_cycloneiii_0_s1_allgrants <= remote_update_cycloneiii_0_s1_grant_vector;
  --remote_update_cycloneiii_0_s1_end_xfer assignment, which is an e_assign
  remote_update_cycloneiii_0_s1_end_xfer <= NOT ((remote_update_cycloneiii_0_s1_waits_for_read OR remote_update_cycloneiii_0_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_remote_update_cycloneiii_0_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_remote_update_cycloneiii_0_s1 <= remote_update_cycloneiii_0_s1_end_xfer AND (((NOT remote_update_cycloneiii_0_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --remote_update_cycloneiii_0_s1_arb_share_counter arbitration counter enable, which is an e_assign
  remote_update_cycloneiii_0_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_remote_update_cycloneiii_0_s1 AND remote_update_cycloneiii_0_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_remote_update_cycloneiii_0_s1 AND NOT remote_update_cycloneiii_0_s1_non_bursting_master_requests));
  --remote_update_cycloneiii_0_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      remote_update_cycloneiii_0_s1_arb_share_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(remote_update_cycloneiii_0_s1_arb_counter_enable) = '1' then 
        remote_update_cycloneiii_0_s1_arb_share_counter <= remote_update_cycloneiii_0_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --remote_update_cycloneiii_0_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      remote_update_cycloneiii_0_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((remote_update_cycloneiii_0_s1_master_qreq_vector AND end_xfer_arb_share_counter_term_remote_update_cycloneiii_0_s1)) OR ((end_xfer_arb_share_counter_term_remote_update_cycloneiii_0_s1 AND NOT remote_update_cycloneiii_0_s1_non_bursting_master_requests)))) = '1' then 
        remote_update_cycloneiii_0_s1_slavearbiterlockenable <= remote_update_cycloneiii_0_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --niosII_openMac_clock_4/out remote_update_cycloneiii_0/s1 arbiterlock, which is an e_assign
  niosII_openMac_clock_4_out_arbiterlock <= remote_update_cycloneiii_0_s1_slavearbiterlockenable AND niosII_openMac_clock_4_out_continuerequest;
  --remote_update_cycloneiii_0_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  remote_update_cycloneiii_0_s1_slavearbiterlockenable2 <= remote_update_cycloneiii_0_s1_arb_share_counter_next_value;
  --niosII_openMac_clock_4/out remote_update_cycloneiii_0/s1 arbiterlock2, which is an e_assign
  niosII_openMac_clock_4_out_arbiterlock2 <= remote_update_cycloneiii_0_s1_slavearbiterlockenable2 AND niosII_openMac_clock_4_out_continuerequest;
  --remote_update_cycloneiii_0_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  remote_update_cycloneiii_0_s1_any_continuerequest <= std_logic'('1');
  --niosII_openMac_clock_4_out_continuerequest continued request, which is an e_assign
  niosII_openMac_clock_4_out_continuerequest <= std_logic'('1');
  internal_niosII_openMac_clock_4_out_qualified_request_remote_update_cycloneiii_0_s1 <= internal_niosII_openMac_clock_4_out_requests_remote_update_cycloneiii_0_s1 AND NOT ((niosII_openMac_clock_4_out_read AND (or_reduce(niosII_openMac_clock_4_out_read_data_valid_remote_update_cycloneiii_0_s1_shift_register))));
  --niosII_openMac_clock_4_out_read_data_valid_remote_update_cycloneiii_0_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  niosII_openMac_clock_4_out_read_data_valid_remote_update_cycloneiii_0_s1_shift_register_in <= ((internal_niosII_openMac_clock_4_out_granted_remote_update_cycloneiii_0_s1 AND niosII_openMac_clock_4_out_read) AND NOT remote_update_cycloneiii_0_s1_waits_for_read) AND NOT (or_reduce(niosII_openMac_clock_4_out_read_data_valid_remote_update_cycloneiii_0_s1_shift_register));
  --shift register p1 niosII_openMac_clock_4_out_read_data_valid_remote_update_cycloneiii_0_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  p1_niosII_openMac_clock_4_out_read_data_valid_remote_update_cycloneiii_0_s1_shift_register <= A_EXT ((niosII_openMac_clock_4_out_read_data_valid_remote_update_cycloneiii_0_s1_shift_register & A_ToStdLogicVector(niosII_openMac_clock_4_out_read_data_valid_remote_update_cycloneiii_0_s1_shift_register_in)), 2);
  --niosII_openMac_clock_4_out_read_data_valid_remote_update_cycloneiii_0_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      niosII_openMac_clock_4_out_read_data_valid_remote_update_cycloneiii_0_s1_shift_register <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      niosII_openMac_clock_4_out_read_data_valid_remote_update_cycloneiii_0_s1_shift_register <= p1_niosII_openMac_clock_4_out_read_data_valid_remote_update_cycloneiii_0_s1_shift_register;
    end if;

  end process;

  --local readdatavalid niosII_openMac_clock_4_out_read_data_valid_remote_update_cycloneiii_0_s1, which is an e_mux
  niosII_openMac_clock_4_out_read_data_valid_remote_update_cycloneiii_0_s1 <= niosII_openMac_clock_4_out_read_data_valid_remote_update_cycloneiii_0_s1_shift_register(1);
  --remote_update_cycloneiii_0_s1_writedata mux, which is an e_mux
  remote_update_cycloneiii_0_s1_writedata <= niosII_openMac_clock_4_out_writedata;
  --master is always granted when requested
  internal_niosII_openMac_clock_4_out_granted_remote_update_cycloneiii_0_s1 <= internal_niosII_openMac_clock_4_out_qualified_request_remote_update_cycloneiii_0_s1;
  --niosII_openMac_clock_4/out saved-grant remote_update_cycloneiii_0/s1, which is an e_assign
  niosII_openMac_clock_4_out_saved_grant_remote_update_cycloneiii_0_s1 <= internal_niosII_openMac_clock_4_out_requests_remote_update_cycloneiii_0_s1;
  --allow new arb cycle for remote_update_cycloneiii_0/s1, which is an e_assign
  remote_update_cycloneiii_0_s1_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  remote_update_cycloneiii_0_s1_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  remote_update_cycloneiii_0_s1_master_qreq_vector <= std_logic'('1');
  --~remote_update_cycloneiii_0_s1_reset assignment, which is an e_assign
  remote_update_cycloneiii_0_s1_reset <= NOT reset_n;
  remote_update_cycloneiii_0_s1_chipselect <= internal_niosII_openMac_clock_4_out_granted_remote_update_cycloneiii_0_s1;
  --remote_update_cycloneiii_0_s1_firsttransfer first transaction, which is an e_assign
  remote_update_cycloneiii_0_s1_firsttransfer <= A_WE_StdLogic((std_logic'(remote_update_cycloneiii_0_s1_begins_xfer) = '1'), remote_update_cycloneiii_0_s1_unreg_firsttransfer, remote_update_cycloneiii_0_s1_reg_firsttransfer);
  --remote_update_cycloneiii_0_s1_unreg_firsttransfer first transaction, which is an e_assign
  remote_update_cycloneiii_0_s1_unreg_firsttransfer <= NOT ((remote_update_cycloneiii_0_s1_slavearbiterlockenable AND remote_update_cycloneiii_0_s1_any_continuerequest));
  --remote_update_cycloneiii_0_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      remote_update_cycloneiii_0_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(remote_update_cycloneiii_0_s1_begins_xfer) = '1' then 
        remote_update_cycloneiii_0_s1_reg_firsttransfer <= remote_update_cycloneiii_0_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --remote_update_cycloneiii_0_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  remote_update_cycloneiii_0_s1_beginbursttransfer_internal <= remote_update_cycloneiii_0_s1_begins_xfer;
  --remote_update_cycloneiii_0_s1_read assignment, which is an e_mux
  remote_update_cycloneiii_0_s1_read <= internal_niosII_openMac_clock_4_out_granted_remote_update_cycloneiii_0_s1 AND niosII_openMac_clock_4_out_read;
  --remote_update_cycloneiii_0_s1_write assignment, which is an e_mux
  remote_update_cycloneiii_0_s1_write <= internal_niosII_openMac_clock_4_out_granted_remote_update_cycloneiii_0_s1 AND niosII_openMac_clock_4_out_write;
  --remote_update_cycloneiii_0_s1_address mux, which is an e_mux
  remote_update_cycloneiii_0_s1_address <= niosII_openMac_clock_4_out_nativeaddress;
  --d1_remote_update_cycloneiii_0_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_remote_update_cycloneiii_0_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_remote_update_cycloneiii_0_s1_end_xfer <= remote_update_cycloneiii_0_s1_end_xfer;
    end if;

  end process;

  --remote_update_cycloneiii_0_s1_waits_for_read in a cycle, which is an e_mux
  remote_update_cycloneiii_0_s1_waits_for_read <= remote_update_cycloneiii_0_s1_in_a_read_cycle AND internal_remote_update_cycloneiii_0_s1_waitrequest_from_sa;
  --remote_update_cycloneiii_0_s1_in_a_read_cycle assignment, which is an e_assign
  remote_update_cycloneiii_0_s1_in_a_read_cycle <= internal_niosII_openMac_clock_4_out_granted_remote_update_cycloneiii_0_s1 AND niosII_openMac_clock_4_out_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= remote_update_cycloneiii_0_s1_in_a_read_cycle;
  --remote_update_cycloneiii_0_s1_waits_for_write in a cycle, which is an e_mux
  remote_update_cycloneiii_0_s1_waits_for_write <= remote_update_cycloneiii_0_s1_in_a_write_cycle AND internal_remote_update_cycloneiii_0_s1_waitrequest_from_sa;
  --remote_update_cycloneiii_0_s1_in_a_write_cycle assignment, which is an e_assign
  remote_update_cycloneiii_0_s1_in_a_write_cycle <= internal_niosII_openMac_clock_4_out_granted_remote_update_cycloneiii_0_s1 AND niosII_openMac_clock_4_out_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= remote_update_cycloneiii_0_s1_in_a_write_cycle;
  wait_for_remote_update_cycloneiii_0_s1_counter <= std_logic'('0');
  --vhdl renameroo for output signals
  niosII_openMac_clock_4_out_granted_remote_update_cycloneiii_0_s1 <= internal_niosII_openMac_clock_4_out_granted_remote_update_cycloneiii_0_s1;
  --vhdl renameroo for output signals
  niosII_openMac_clock_4_out_qualified_request_remote_update_cycloneiii_0_s1 <= internal_niosII_openMac_clock_4_out_qualified_request_remote_update_cycloneiii_0_s1;
  --vhdl renameroo for output signals
  niosII_openMac_clock_4_out_requests_remote_update_cycloneiii_0_s1 <= internal_niosII_openMac_clock_4_out_requests_remote_update_cycloneiii_0_s1;
  --vhdl renameroo for output signals
  remote_update_cycloneiii_0_s1_waitrequest_from_sa <= internal_remote_update_cycloneiii_0_s1_waitrequest_from_sa;
--synthesis translate_off
    --remote_update_cycloneiii_0/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity rdv_fifo_for_ap_cpu_data_master_to_sdram_0_s1_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC;
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity rdv_fifo_for_ap_cpu_data_master_to_sdram_0_s1_module;


architecture europa of rdv_fifo_for_ap_cpu_data_master_to_sdram_0_s1_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal full_3 :  STD_LOGIC;
                signal full_4 :  STD_LOGIC;
                signal full_5 :  STD_LOGIC;
                signal full_6 :  STD_LOGIC;
                signal full_7 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC;
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC;
                signal p2_full_2 :  STD_LOGIC;
                signal p2_stage_2 :  STD_LOGIC;
                signal p3_full_3 :  STD_LOGIC;
                signal p3_stage_3 :  STD_LOGIC;
                signal p4_full_4 :  STD_LOGIC;
                signal p4_stage_4 :  STD_LOGIC;
                signal p5_full_5 :  STD_LOGIC;
                signal p5_stage_5 :  STD_LOGIC;
                signal p6_full_6 :  STD_LOGIC;
                signal p6_stage_6 :  STD_LOGIC;
                signal stage_0 :  STD_LOGIC;
                signal stage_1 :  STD_LOGIC;
                signal stage_2 :  STD_LOGIC;
                signal stage_3 :  STD_LOGIC;
                signal stage_4 :  STD_LOGIC;
                signal stage_5 :  STD_LOGIC;
                signal stage_6 :  STD_LOGIC;
                signal updated_one_count :  STD_LOGIC_VECTOR (3 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_6;
  empty <= NOT(full_0);
  full_7 <= std_logic'('0');
  --data_6, which is an e_mux
  p6_stage_6 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_7 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_6 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_6))))) = '1' then 
        if std_logic'(((sync_reset AND full_6) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_7))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_6 <= std_logic'('0');
        else
          stage_6 <= p6_stage_6;
        end if;
      end if;
    end if;

  end process;

  --control_6, which is an e_mux
  p6_full_6 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_5))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_6 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_6 <= std_logic'('0');
        else
          full_6 <= p6_full_6;
        end if;
      end if;
    end if;

  end process;

  --data_5, which is an e_mux
  p5_stage_5 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_6 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_6);
  --data_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_5))))) = '1' then 
        if std_logic'(((sync_reset AND full_5) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_6))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_5 <= std_logic'('0');
        else
          stage_5 <= p5_stage_5;
        end if;
      end if;
    end if;

  end process;

  --control_5, which is an e_mux
  p5_full_5 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_4, full_6);
  --control_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_5 <= std_logic'('0');
        else
          full_5 <= p5_full_5;
        end if;
      end if;
    end if;

  end process;

  --data_4, which is an e_mux
  p4_stage_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_5 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_5);
  --data_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_4))))) = '1' then 
        if std_logic'(((sync_reset AND full_4) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_5))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_4 <= std_logic'('0');
        else
          stage_4 <= p4_stage_4;
        end if;
      end if;
    end if;

  end process;

  --control_4, which is an e_mux
  p4_full_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_3, full_5);
  --control_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_4 <= std_logic'('0');
        else
          full_4 <= p4_full_4;
        end if;
      end if;
    end if;

  end process;

  --data_3, which is an e_mux
  p3_stage_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_4 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_4);
  --data_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_3))))) = '1' then 
        if std_logic'(((sync_reset AND full_3) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_4))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_3 <= std_logic'('0');
        else
          stage_3 <= p3_stage_3;
        end if;
      end if;
    end if;

  end process;

  --control_3, which is an e_mux
  p3_full_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_2, full_4);
  --control_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_3 <= std_logic'('0');
        else
          full_3 <= p3_full_3;
        end if;
      end if;
    end if;

  end process;

  --data_2, which is an e_mux
  p2_stage_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_3 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_3);
  --data_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_2))))) = '1' then 
        if std_logic'(((sync_reset AND full_2) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_3))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_2 <= std_logic'('0');
        else
          stage_2 <= p2_stage_2;
        end if;
      end if;
    end if;

  end process;

  --control_2, which is an e_mux
  p2_full_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_1, full_3);
  --control_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_2 <= std_logic'('0');
        else
          full_2 <= p2_full_2;
        end if;
      end if;
    end if;

  end process;

  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_2);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic'('0');
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_0, full_2);
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic'('0');
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 4);
  one_count_minus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 4);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("000") & (A_TOSTDLOGICVECTOR(data_in))), A_WE_StdLogicVector((std_logic'(((((read AND (data_in)) AND write) AND (stage_0)))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (data_in)))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (stage_0)))) = '1'), one_count_minus_one, how_many_ones))))))), 4);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity rdv_fifo_for_ap_cpu_instruction_master_to_sdram_0_s1_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC;
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity rdv_fifo_for_ap_cpu_instruction_master_to_sdram_0_s1_module;


architecture europa of rdv_fifo_for_ap_cpu_instruction_master_to_sdram_0_s1_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal full_3 :  STD_LOGIC;
                signal full_4 :  STD_LOGIC;
                signal full_5 :  STD_LOGIC;
                signal full_6 :  STD_LOGIC;
                signal full_7 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC;
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC;
                signal p2_full_2 :  STD_LOGIC;
                signal p2_stage_2 :  STD_LOGIC;
                signal p3_full_3 :  STD_LOGIC;
                signal p3_stage_3 :  STD_LOGIC;
                signal p4_full_4 :  STD_LOGIC;
                signal p4_stage_4 :  STD_LOGIC;
                signal p5_full_5 :  STD_LOGIC;
                signal p5_stage_5 :  STD_LOGIC;
                signal p6_full_6 :  STD_LOGIC;
                signal p6_stage_6 :  STD_LOGIC;
                signal stage_0 :  STD_LOGIC;
                signal stage_1 :  STD_LOGIC;
                signal stage_2 :  STD_LOGIC;
                signal stage_3 :  STD_LOGIC;
                signal stage_4 :  STD_LOGIC;
                signal stage_5 :  STD_LOGIC;
                signal stage_6 :  STD_LOGIC;
                signal updated_one_count :  STD_LOGIC_VECTOR (3 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_6;
  empty <= NOT(full_0);
  full_7 <= std_logic'('0');
  --data_6, which is an e_mux
  p6_stage_6 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_7 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_6 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_6))))) = '1' then 
        if std_logic'(((sync_reset AND full_6) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_7))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_6 <= std_logic'('0');
        else
          stage_6 <= p6_stage_6;
        end if;
      end if;
    end if;

  end process;

  --control_6, which is an e_mux
  p6_full_6 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_5))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_6 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_6 <= std_logic'('0');
        else
          full_6 <= p6_full_6;
        end if;
      end if;
    end if;

  end process;

  --data_5, which is an e_mux
  p5_stage_5 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_6 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_6);
  --data_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_5))))) = '1' then 
        if std_logic'(((sync_reset AND full_5) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_6))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_5 <= std_logic'('0');
        else
          stage_5 <= p5_stage_5;
        end if;
      end if;
    end if;

  end process;

  --control_5, which is an e_mux
  p5_full_5 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_4, full_6);
  --control_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_5 <= std_logic'('0');
        else
          full_5 <= p5_full_5;
        end if;
      end if;
    end if;

  end process;

  --data_4, which is an e_mux
  p4_stage_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_5 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_5);
  --data_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_4))))) = '1' then 
        if std_logic'(((sync_reset AND full_4) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_5))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_4 <= std_logic'('0');
        else
          stage_4 <= p4_stage_4;
        end if;
      end if;
    end if;

  end process;

  --control_4, which is an e_mux
  p4_full_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_3, full_5);
  --control_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_4 <= std_logic'('0');
        else
          full_4 <= p4_full_4;
        end if;
      end if;
    end if;

  end process;

  --data_3, which is an e_mux
  p3_stage_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_4 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_4);
  --data_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_3))))) = '1' then 
        if std_logic'(((sync_reset AND full_3) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_4))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_3 <= std_logic'('0');
        else
          stage_3 <= p3_stage_3;
        end if;
      end if;
    end if;

  end process;

  --control_3, which is an e_mux
  p3_full_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_2, full_4);
  --control_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_3 <= std_logic'('0');
        else
          full_3 <= p3_full_3;
        end if;
      end if;
    end if;

  end process;

  --data_2, which is an e_mux
  p2_stage_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_3 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_3);
  --data_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_2))))) = '1' then 
        if std_logic'(((sync_reset AND full_2) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_3))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_2 <= std_logic'('0');
        else
          stage_2 <= p2_stage_2;
        end if;
      end if;
    end if;

  end process;

  --control_2, which is an e_mux
  p2_full_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_1, full_3);
  --control_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_2 <= std_logic'('0');
        else
          full_2 <= p2_full_2;
        end if;
      end if;
    end if;

  end process;

  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_2);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic'('0');
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_0, full_2);
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic'('0');
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 4);
  one_count_minus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 4);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("000") & (A_TOSTDLOGICVECTOR(data_in))), A_WE_StdLogicVector((std_logic'(((((read AND (data_in)) AND write) AND (stage_0)))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (data_in)))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (stage_0)))) = '1'), one_count_minus_one, how_many_ones))))))), 4);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity sdram_0_s1_arbitrator is 
        port (
              -- inputs:
                 signal ap_cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (25 DOWNTO 0);
                 signal ap_cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal ap_cpu_data_master_read : IN STD_LOGIC;
                 signal ap_cpu_data_master_waitrequest : IN STD_LOGIC;
                 signal ap_cpu_data_master_write : IN STD_LOGIC;
                 signal ap_cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal ap_cpu_instruction_master_address_to_slave : IN STD_LOGIC_VECTOR (25 DOWNTO 0);
                 signal ap_cpu_instruction_master_latency_counter : IN STD_LOGIC;
                 signal ap_cpu_instruction_master_read : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sdram_0_s1_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal sdram_0_s1_readdatavalid : IN STD_LOGIC;
                 signal sdram_0_s1_waitrequest : IN STD_LOGIC;

              -- outputs:
                 signal ap_cpu_data_master_granted_sdram_0_s1 : OUT STD_LOGIC;
                 signal ap_cpu_data_master_qualified_request_sdram_0_s1 : OUT STD_LOGIC;
                 signal ap_cpu_data_master_read_data_valid_sdram_0_s1 : OUT STD_LOGIC;
                 signal ap_cpu_data_master_read_data_valid_sdram_0_s1_shift_register : OUT STD_LOGIC;
                 signal ap_cpu_data_master_requests_sdram_0_s1 : OUT STD_LOGIC;
                 signal ap_cpu_instruction_master_granted_sdram_0_s1 : OUT STD_LOGIC;
                 signal ap_cpu_instruction_master_qualified_request_sdram_0_s1 : OUT STD_LOGIC;
                 signal ap_cpu_instruction_master_read_data_valid_sdram_0_s1 : OUT STD_LOGIC;
                 signal ap_cpu_instruction_master_read_data_valid_sdram_0_s1_shift_register : OUT STD_LOGIC;
                 signal ap_cpu_instruction_master_requests_sdram_0_s1 : OUT STD_LOGIC;
                 signal d1_sdram_0_s1_end_xfer : OUT STD_LOGIC;
                 signal sdram_0_s1_address : OUT STD_LOGIC_VECTOR (21 DOWNTO 0);
                 signal sdram_0_s1_byteenable_n : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal sdram_0_s1_chipselect : OUT STD_LOGIC;
                 signal sdram_0_s1_read_n : OUT STD_LOGIC;
                 signal sdram_0_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal sdram_0_s1_reset_n : OUT STD_LOGIC;
                 signal sdram_0_s1_waitrequest_from_sa : OUT STD_LOGIC;
                 signal sdram_0_s1_write_n : OUT STD_LOGIC;
                 signal sdram_0_s1_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
              );
end entity sdram_0_s1_arbitrator;


architecture europa of sdram_0_s1_arbitrator is
component rdv_fifo_for_ap_cpu_data_master_to_sdram_0_s1_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC;
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component rdv_fifo_for_ap_cpu_data_master_to_sdram_0_s1_module;

component rdv_fifo_for_ap_cpu_instruction_master_to_sdram_0_s1_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC;
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component rdv_fifo_for_ap_cpu_instruction_master_to_sdram_0_s1_module;

                signal ap_cpu_data_master_arbiterlock :  STD_LOGIC;
                signal ap_cpu_data_master_arbiterlock2 :  STD_LOGIC;
                signal ap_cpu_data_master_continuerequest :  STD_LOGIC;
                signal ap_cpu_data_master_rdv_fifo_empty_sdram_0_s1 :  STD_LOGIC;
                signal ap_cpu_data_master_rdv_fifo_output_from_sdram_0_s1 :  STD_LOGIC;
                signal ap_cpu_data_master_saved_grant_sdram_0_s1 :  STD_LOGIC;
                signal ap_cpu_instruction_master_arbiterlock :  STD_LOGIC;
                signal ap_cpu_instruction_master_arbiterlock2 :  STD_LOGIC;
                signal ap_cpu_instruction_master_continuerequest :  STD_LOGIC;
                signal ap_cpu_instruction_master_rdv_fifo_empty_sdram_0_s1 :  STD_LOGIC;
                signal ap_cpu_instruction_master_rdv_fifo_output_from_sdram_0_s1 :  STD_LOGIC;
                signal ap_cpu_instruction_master_saved_grant_sdram_0_s1 :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_sdram_0_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_ap_cpu_data_master_granted_sdram_0_s1 :  STD_LOGIC;
                signal internal_ap_cpu_data_master_qualified_request_sdram_0_s1 :  STD_LOGIC;
                signal internal_ap_cpu_data_master_read_data_valid_sdram_0_s1_shift_register :  STD_LOGIC;
                signal internal_ap_cpu_data_master_requests_sdram_0_s1 :  STD_LOGIC;
                signal internal_ap_cpu_instruction_master_granted_sdram_0_s1 :  STD_LOGIC;
                signal internal_ap_cpu_instruction_master_qualified_request_sdram_0_s1 :  STD_LOGIC;
                signal internal_ap_cpu_instruction_master_requests_sdram_0_s1 :  STD_LOGIC;
                signal internal_sdram_0_s1_waitrequest_from_sa :  STD_LOGIC;
                signal last_cycle_ap_cpu_data_master_granted_slave_sdram_0_s1 :  STD_LOGIC;
                signal last_cycle_ap_cpu_instruction_master_granted_slave_sdram_0_s1 :  STD_LOGIC;
                signal module_input10 :  STD_LOGIC;
                signal module_input11 :  STD_LOGIC;
                signal module_input6 :  STD_LOGIC;
                signal module_input7 :  STD_LOGIC;
                signal module_input8 :  STD_LOGIC;
                signal module_input9 :  STD_LOGIC;
                signal sdram_0_s1_allgrants :  STD_LOGIC;
                signal sdram_0_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal sdram_0_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal sdram_0_s1_any_continuerequest :  STD_LOGIC;
                signal sdram_0_s1_arb_addend :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal sdram_0_s1_arb_counter_enable :  STD_LOGIC;
                signal sdram_0_s1_arb_share_counter :  STD_LOGIC;
                signal sdram_0_s1_arb_share_counter_next_value :  STD_LOGIC;
                signal sdram_0_s1_arb_share_set_values :  STD_LOGIC;
                signal sdram_0_s1_arb_winner :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal sdram_0_s1_arbitration_holdoff_internal :  STD_LOGIC;
                signal sdram_0_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal sdram_0_s1_begins_xfer :  STD_LOGIC;
                signal sdram_0_s1_chosen_master_double_vector :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal sdram_0_s1_chosen_master_rot_left :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal sdram_0_s1_end_xfer :  STD_LOGIC;
                signal sdram_0_s1_firsttransfer :  STD_LOGIC;
                signal sdram_0_s1_grant_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal sdram_0_s1_in_a_read_cycle :  STD_LOGIC;
                signal sdram_0_s1_in_a_write_cycle :  STD_LOGIC;
                signal sdram_0_s1_master_qreq_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal sdram_0_s1_move_on_to_next_transaction :  STD_LOGIC;
                signal sdram_0_s1_non_bursting_master_requests :  STD_LOGIC;
                signal sdram_0_s1_readdatavalid_from_sa :  STD_LOGIC;
                signal sdram_0_s1_reg_firsttransfer :  STD_LOGIC;
                signal sdram_0_s1_saved_chosen_master_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal sdram_0_s1_slavearbiterlockenable :  STD_LOGIC;
                signal sdram_0_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal sdram_0_s1_unreg_firsttransfer :  STD_LOGIC;
                signal sdram_0_s1_waits_for_read :  STD_LOGIC;
                signal sdram_0_s1_waits_for_write :  STD_LOGIC;
                signal shifted_address_to_sdram_0_s1_from_ap_cpu_data_master :  STD_LOGIC_VECTOR (25 DOWNTO 0);
                signal shifted_address_to_sdram_0_s1_from_ap_cpu_instruction_master :  STD_LOGIC_VECTOR (25 DOWNTO 0);
                signal wait_for_sdram_0_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT sdram_0_s1_end_xfer;
    end if;

  end process;

  sdram_0_s1_begins_xfer <= NOT d1_reasons_to_wait AND ((internal_ap_cpu_data_master_qualified_request_sdram_0_s1 OR internal_ap_cpu_instruction_master_qualified_request_sdram_0_s1));
  --assign sdram_0_s1_readdatavalid_from_sa = sdram_0_s1_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  sdram_0_s1_readdatavalid_from_sa <= sdram_0_s1_readdatavalid;
  --assign sdram_0_s1_readdata_from_sa = sdram_0_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  sdram_0_s1_readdata_from_sa <= sdram_0_s1_readdata;
  internal_ap_cpu_data_master_requests_sdram_0_s1 <= to_std_logic(((Std_Logic_Vector'(ap_cpu_data_master_address_to_slave(25 DOWNTO 24) & std_logic_vector'("000000000000000000000000")) = std_logic_vector'("10000000000000000000000000")))) AND ((ap_cpu_data_master_read OR ap_cpu_data_master_write));
  --assign sdram_0_s1_waitrequest_from_sa = sdram_0_s1_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_sdram_0_s1_waitrequest_from_sa <= sdram_0_s1_waitrequest;
  --sdram_0_s1_arb_share_counter set values, which is an e_mux
  sdram_0_s1_arb_share_set_values <= std_logic'('1');
  --sdram_0_s1_non_bursting_master_requests mux, which is an e_mux
  sdram_0_s1_non_bursting_master_requests <= ((internal_ap_cpu_data_master_requests_sdram_0_s1 OR internal_ap_cpu_instruction_master_requests_sdram_0_s1) OR internal_ap_cpu_data_master_requests_sdram_0_s1) OR internal_ap_cpu_instruction_master_requests_sdram_0_s1;
  --sdram_0_s1_any_bursting_master_saved_grant mux, which is an e_mux
  sdram_0_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --sdram_0_s1_arb_share_counter_next_value assignment, which is an e_assign
  sdram_0_s1_arb_share_counter_next_value <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(sdram_0_s1_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(sdram_0_s1_arb_share_set_values))) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(sdram_0_s1_arb_share_counter) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(sdram_0_s1_arb_share_counter))) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))));
  --sdram_0_s1_allgrants all slave grants, which is an e_mux
  sdram_0_s1_allgrants <= (((or_reduce(sdram_0_s1_grant_vector)) OR (or_reduce(sdram_0_s1_grant_vector))) OR (or_reduce(sdram_0_s1_grant_vector))) OR (or_reduce(sdram_0_s1_grant_vector));
  --sdram_0_s1_end_xfer assignment, which is an e_assign
  sdram_0_s1_end_xfer <= NOT ((sdram_0_s1_waits_for_read OR sdram_0_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_sdram_0_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_sdram_0_s1 <= sdram_0_s1_end_xfer AND (((NOT sdram_0_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --sdram_0_s1_arb_share_counter arbitration counter enable, which is an e_assign
  sdram_0_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_sdram_0_s1 AND sdram_0_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_sdram_0_s1 AND NOT sdram_0_s1_non_bursting_master_requests));
  --sdram_0_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sdram_0_s1_arb_share_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(sdram_0_s1_arb_counter_enable) = '1' then 
        sdram_0_s1_arb_share_counter <= sdram_0_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --sdram_0_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sdram_0_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((or_reduce(sdram_0_s1_master_qreq_vector) AND end_xfer_arb_share_counter_term_sdram_0_s1)) OR ((end_xfer_arb_share_counter_term_sdram_0_s1 AND NOT sdram_0_s1_non_bursting_master_requests)))) = '1' then 
        sdram_0_s1_slavearbiterlockenable <= sdram_0_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --ap_cpu/data_master sdram_0/s1 arbiterlock, which is an e_assign
  ap_cpu_data_master_arbiterlock <= sdram_0_s1_slavearbiterlockenable AND ap_cpu_data_master_continuerequest;
  --sdram_0_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  sdram_0_s1_slavearbiterlockenable2 <= sdram_0_s1_arb_share_counter_next_value;
  --ap_cpu/data_master sdram_0/s1 arbiterlock2, which is an e_assign
  ap_cpu_data_master_arbiterlock2 <= sdram_0_s1_slavearbiterlockenable2 AND ap_cpu_data_master_continuerequest;
  --ap_cpu/instruction_master sdram_0/s1 arbiterlock, which is an e_assign
  ap_cpu_instruction_master_arbiterlock <= sdram_0_s1_slavearbiterlockenable AND ap_cpu_instruction_master_continuerequest;
  --ap_cpu/instruction_master sdram_0/s1 arbiterlock2, which is an e_assign
  ap_cpu_instruction_master_arbiterlock2 <= sdram_0_s1_slavearbiterlockenable2 AND ap_cpu_instruction_master_continuerequest;
  --ap_cpu/instruction_master granted sdram_0/s1 last time, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      last_cycle_ap_cpu_instruction_master_granted_slave_sdram_0_s1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      last_cycle_ap_cpu_instruction_master_granted_slave_sdram_0_s1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(ap_cpu_instruction_master_saved_grant_sdram_0_s1) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((sdram_0_s1_arbitration_holdoff_internal OR NOT internal_ap_cpu_instruction_master_requests_sdram_0_s1))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_ap_cpu_instruction_master_granted_slave_sdram_0_s1))))));
    end if;

  end process;

  --ap_cpu_instruction_master_continuerequest continued request, which is an e_mux
  ap_cpu_instruction_master_continuerequest <= last_cycle_ap_cpu_instruction_master_granted_slave_sdram_0_s1 AND internal_ap_cpu_instruction_master_requests_sdram_0_s1;
  --sdram_0_s1_any_continuerequest at least one master continues requesting, which is an e_mux
  sdram_0_s1_any_continuerequest <= ap_cpu_instruction_master_continuerequest OR ap_cpu_data_master_continuerequest;
  internal_ap_cpu_data_master_qualified_request_sdram_0_s1 <= internal_ap_cpu_data_master_requests_sdram_0_s1 AND NOT (((((ap_cpu_data_master_read AND ((NOT ap_cpu_data_master_waitrequest OR (internal_ap_cpu_data_master_read_data_valid_sdram_0_s1_shift_register))))) OR (((NOT ap_cpu_data_master_waitrequest) AND ap_cpu_data_master_write))) OR ap_cpu_instruction_master_arbiterlock));
  --unique name for sdram_0_s1_move_on_to_next_transaction, which is an e_assign
  sdram_0_s1_move_on_to_next_transaction <= sdram_0_s1_readdatavalid_from_sa;
  --rdv_fifo_for_ap_cpu_data_master_to_sdram_0_s1, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_ap_cpu_data_master_to_sdram_0_s1 : rdv_fifo_for_ap_cpu_data_master_to_sdram_0_s1_module
    port map(
      data_out => ap_cpu_data_master_rdv_fifo_output_from_sdram_0_s1,
      empty => open,
      fifo_contains_ones_n => ap_cpu_data_master_rdv_fifo_empty_sdram_0_s1,
      full => open,
      clear_fifo => module_input6,
      clk => clk,
      data_in => internal_ap_cpu_data_master_granted_sdram_0_s1,
      read => sdram_0_s1_move_on_to_next_transaction,
      reset_n => reset_n,
      sync_reset => module_input7,
      write => module_input8
    );

  module_input6 <= std_logic'('0');
  module_input7 <= std_logic'('0');
  module_input8 <= in_a_read_cycle AND NOT sdram_0_s1_waits_for_read;

  internal_ap_cpu_data_master_read_data_valid_sdram_0_s1_shift_register <= NOT ap_cpu_data_master_rdv_fifo_empty_sdram_0_s1;
  --local readdatavalid ap_cpu_data_master_read_data_valid_sdram_0_s1, which is an e_mux
  ap_cpu_data_master_read_data_valid_sdram_0_s1 <= ((sdram_0_s1_readdatavalid_from_sa AND ap_cpu_data_master_rdv_fifo_output_from_sdram_0_s1)) AND NOT ap_cpu_data_master_rdv_fifo_empty_sdram_0_s1;
  --sdram_0_s1_writedata mux, which is an e_mux
  sdram_0_s1_writedata <= ap_cpu_data_master_writedata;
  internal_ap_cpu_instruction_master_requests_sdram_0_s1 <= ((to_std_logic(((Std_Logic_Vector'(ap_cpu_instruction_master_address_to_slave(25 DOWNTO 24) & std_logic_vector'("000000000000000000000000")) = std_logic_vector'("10000000000000000000000000")))) AND (ap_cpu_instruction_master_read))) AND ap_cpu_instruction_master_read;
  --ap_cpu/data_master granted sdram_0/s1 last time, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      last_cycle_ap_cpu_data_master_granted_slave_sdram_0_s1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      last_cycle_ap_cpu_data_master_granted_slave_sdram_0_s1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(ap_cpu_data_master_saved_grant_sdram_0_s1) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((sdram_0_s1_arbitration_holdoff_internal OR NOT internal_ap_cpu_data_master_requests_sdram_0_s1))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_ap_cpu_data_master_granted_slave_sdram_0_s1))))));
    end if;

  end process;

  --ap_cpu_data_master_continuerequest continued request, which is an e_mux
  ap_cpu_data_master_continuerequest <= last_cycle_ap_cpu_data_master_granted_slave_sdram_0_s1 AND internal_ap_cpu_data_master_requests_sdram_0_s1;
  internal_ap_cpu_instruction_master_qualified_request_sdram_0_s1 <= internal_ap_cpu_instruction_master_requests_sdram_0_s1 AND NOT ((((ap_cpu_instruction_master_read AND to_std_logic((((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(ap_cpu_instruction_master_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))) OR ((std_logic_vector'("00000000000000000000000000000001")<(std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(ap_cpu_instruction_master_latency_counter)))))))))) OR ap_cpu_data_master_arbiterlock));
  --rdv_fifo_for_ap_cpu_instruction_master_to_sdram_0_s1, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_ap_cpu_instruction_master_to_sdram_0_s1 : rdv_fifo_for_ap_cpu_instruction_master_to_sdram_0_s1_module
    port map(
      data_out => ap_cpu_instruction_master_rdv_fifo_output_from_sdram_0_s1,
      empty => open,
      fifo_contains_ones_n => ap_cpu_instruction_master_rdv_fifo_empty_sdram_0_s1,
      full => open,
      clear_fifo => module_input9,
      clk => clk,
      data_in => internal_ap_cpu_instruction_master_granted_sdram_0_s1,
      read => sdram_0_s1_move_on_to_next_transaction,
      reset_n => reset_n,
      sync_reset => module_input10,
      write => module_input11
    );

  module_input9 <= std_logic'('0');
  module_input10 <= std_logic'('0');
  module_input11 <= in_a_read_cycle AND NOT sdram_0_s1_waits_for_read;

  ap_cpu_instruction_master_read_data_valid_sdram_0_s1_shift_register <= NOT ap_cpu_instruction_master_rdv_fifo_empty_sdram_0_s1;
  --local readdatavalid ap_cpu_instruction_master_read_data_valid_sdram_0_s1, which is an e_mux
  ap_cpu_instruction_master_read_data_valid_sdram_0_s1 <= ((sdram_0_s1_readdatavalid_from_sa AND ap_cpu_instruction_master_rdv_fifo_output_from_sdram_0_s1)) AND NOT ap_cpu_instruction_master_rdv_fifo_empty_sdram_0_s1;
  --allow new arb cycle for sdram_0/s1, which is an e_assign
  sdram_0_s1_allow_new_arb_cycle <= NOT ap_cpu_data_master_arbiterlock AND NOT ap_cpu_instruction_master_arbiterlock;
  --ap_cpu/instruction_master assignment into master qualified-requests vector for sdram_0/s1, which is an e_assign
  sdram_0_s1_master_qreq_vector(0) <= internal_ap_cpu_instruction_master_qualified_request_sdram_0_s1;
  --ap_cpu/instruction_master grant sdram_0/s1, which is an e_assign
  internal_ap_cpu_instruction_master_granted_sdram_0_s1 <= sdram_0_s1_grant_vector(0);
  --ap_cpu/instruction_master saved-grant sdram_0/s1, which is an e_assign
  ap_cpu_instruction_master_saved_grant_sdram_0_s1 <= sdram_0_s1_arb_winner(0) AND internal_ap_cpu_instruction_master_requests_sdram_0_s1;
  --ap_cpu/data_master assignment into master qualified-requests vector for sdram_0/s1, which is an e_assign
  sdram_0_s1_master_qreq_vector(1) <= internal_ap_cpu_data_master_qualified_request_sdram_0_s1;
  --ap_cpu/data_master grant sdram_0/s1, which is an e_assign
  internal_ap_cpu_data_master_granted_sdram_0_s1 <= sdram_0_s1_grant_vector(1);
  --ap_cpu/data_master saved-grant sdram_0/s1, which is an e_assign
  ap_cpu_data_master_saved_grant_sdram_0_s1 <= sdram_0_s1_arb_winner(1) AND internal_ap_cpu_data_master_requests_sdram_0_s1;
  --sdram_0/s1 chosen-master double-vector, which is an e_assign
  sdram_0_s1_chosen_master_double_vector <= A_EXT (((std_logic_vector'("0") & ((sdram_0_s1_master_qreq_vector & sdram_0_s1_master_qreq_vector))) AND (((std_logic_vector'("0") & (Std_Logic_Vector'(NOT sdram_0_s1_master_qreq_vector & NOT sdram_0_s1_master_qreq_vector))) + (std_logic_vector'("000") & (sdram_0_s1_arb_addend))))), 4);
  --stable onehot encoding of arb winner
  sdram_0_s1_arb_winner <= A_WE_StdLogicVector((std_logic'(((sdram_0_s1_allow_new_arb_cycle AND or_reduce(sdram_0_s1_grant_vector)))) = '1'), sdram_0_s1_grant_vector, sdram_0_s1_saved_chosen_master_vector);
  --saved sdram_0_s1_grant_vector, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sdram_0_s1_saved_chosen_master_vector <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      if std_logic'(sdram_0_s1_allow_new_arb_cycle) = '1' then 
        sdram_0_s1_saved_chosen_master_vector <= A_WE_StdLogicVector((std_logic'(or_reduce(sdram_0_s1_grant_vector)) = '1'), sdram_0_s1_grant_vector, sdram_0_s1_saved_chosen_master_vector);
      end if;
    end if;

  end process;

  --onehot encoding of chosen master
  sdram_0_s1_grant_vector <= Std_Logic_Vector'(A_ToStdLogicVector(((sdram_0_s1_chosen_master_double_vector(1) OR sdram_0_s1_chosen_master_double_vector(3)))) & A_ToStdLogicVector(((sdram_0_s1_chosen_master_double_vector(0) OR sdram_0_s1_chosen_master_double_vector(2)))));
  --sdram_0/s1 chosen master rotated left, which is an e_assign
  sdram_0_s1_chosen_master_rot_left <= A_EXT (A_WE_StdLogicVector((((A_SLL(sdram_0_s1_arb_winner,std_logic_vector'("00000000000000000000000000000001")))) /= std_logic_vector'("00")), (std_logic_vector'("000000000000000000000000000000") & ((A_SLL(sdram_0_s1_arb_winner,std_logic_vector'("00000000000000000000000000000001"))))), std_logic_vector'("00000000000000000000000000000001")), 2);
  --sdram_0/s1's addend for next-master-grant
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sdram_0_s1_arb_addend <= std_logic_vector'("01");
    elsif clk'event and clk = '1' then
      if std_logic'(or_reduce(sdram_0_s1_grant_vector)) = '1' then 
        sdram_0_s1_arb_addend <= A_WE_StdLogicVector((std_logic'(sdram_0_s1_end_xfer) = '1'), sdram_0_s1_chosen_master_rot_left, sdram_0_s1_grant_vector);
      end if;
    end if;

  end process;

  --sdram_0_s1_reset_n assignment, which is an e_assign
  sdram_0_s1_reset_n <= reset_n;
  sdram_0_s1_chipselect <= internal_ap_cpu_data_master_granted_sdram_0_s1 OR internal_ap_cpu_instruction_master_granted_sdram_0_s1;
  --sdram_0_s1_firsttransfer first transaction, which is an e_assign
  sdram_0_s1_firsttransfer <= A_WE_StdLogic((std_logic'(sdram_0_s1_begins_xfer) = '1'), sdram_0_s1_unreg_firsttransfer, sdram_0_s1_reg_firsttransfer);
  --sdram_0_s1_unreg_firsttransfer first transaction, which is an e_assign
  sdram_0_s1_unreg_firsttransfer <= NOT ((sdram_0_s1_slavearbiterlockenable AND sdram_0_s1_any_continuerequest));
  --sdram_0_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sdram_0_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(sdram_0_s1_begins_xfer) = '1' then 
        sdram_0_s1_reg_firsttransfer <= sdram_0_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --sdram_0_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  sdram_0_s1_beginbursttransfer_internal <= sdram_0_s1_begins_xfer;
  --sdram_0_s1_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  sdram_0_s1_arbitration_holdoff_internal <= sdram_0_s1_begins_xfer AND sdram_0_s1_firsttransfer;
  --~sdram_0_s1_read_n assignment, which is an e_mux
  sdram_0_s1_read_n <= NOT ((((internal_ap_cpu_data_master_granted_sdram_0_s1 AND ap_cpu_data_master_read)) OR ((internal_ap_cpu_instruction_master_granted_sdram_0_s1 AND ap_cpu_instruction_master_read))));
  --~sdram_0_s1_write_n assignment, which is an e_mux
  sdram_0_s1_write_n <= NOT ((internal_ap_cpu_data_master_granted_sdram_0_s1 AND ap_cpu_data_master_write));
  shifted_address_to_sdram_0_s1_from_ap_cpu_data_master <= ap_cpu_data_master_address_to_slave;
  --sdram_0_s1_address mux, which is an e_mux
  sdram_0_s1_address <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_ap_cpu_data_master_granted_sdram_0_s1)) = '1'), (A_SRL(shifted_address_to_sdram_0_s1_from_ap_cpu_data_master,std_logic_vector'("00000000000000000000000000000010"))), (A_SRL(shifted_address_to_sdram_0_s1_from_ap_cpu_instruction_master,std_logic_vector'("00000000000000000000000000000010")))), 22);
  shifted_address_to_sdram_0_s1_from_ap_cpu_instruction_master <= ap_cpu_instruction_master_address_to_slave;
  --d1_sdram_0_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_sdram_0_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_sdram_0_s1_end_xfer <= sdram_0_s1_end_xfer;
    end if;

  end process;

  --sdram_0_s1_waits_for_read in a cycle, which is an e_mux
  sdram_0_s1_waits_for_read <= sdram_0_s1_in_a_read_cycle AND internal_sdram_0_s1_waitrequest_from_sa;
  --sdram_0_s1_in_a_read_cycle assignment, which is an e_assign
  sdram_0_s1_in_a_read_cycle <= ((internal_ap_cpu_data_master_granted_sdram_0_s1 AND ap_cpu_data_master_read)) OR ((internal_ap_cpu_instruction_master_granted_sdram_0_s1 AND ap_cpu_instruction_master_read));
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= sdram_0_s1_in_a_read_cycle;
  --sdram_0_s1_waits_for_write in a cycle, which is an e_mux
  sdram_0_s1_waits_for_write <= sdram_0_s1_in_a_write_cycle AND internal_sdram_0_s1_waitrequest_from_sa;
  --sdram_0_s1_in_a_write_cycle assignment, which is an e_assign
  sdram_0_s1_in_a_write_cycle <= internal_ap_cpu_data_master_granted_sdram_0_s1 AND ap_cpu_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= sdram_0_s1_in_a_write_cycle;
  wait_for_sdram_0_s1_counter <= std_logic'('0');
  --~sdram_0_s1_byteenable_n byte enable port mux, which is an e_mux
  sdram_0_s1_byteenable_n <= A_EXT (NOT (A_WE_StdLogicVector((std_logic'((internal_ap_cpu_data_master_granted_sdram_0_s1)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (ap_cpu_data_master_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001")))), 4);
  --vhdl renameroo for output signals
  ap_cpu_data_master_granted_sdram_0_s1 <= internal_ap_cpu_data_master_granted_sdram_0_s1;
  --vhdl renameroo for output signals
  ap_cpu_data_master_qualified_request_sdram_0_s1 <= internal_ap_cpu_data_master_qualified_request_sdram_0_s1;
  --vhdl renameroo for output signals
  ap_cpu_data_master_read_data_valid_sdram_0_s1_shift_register <= internal_ap_cpu_data_master_read_data_valid_sdram_0_s1_shift_register;
  --vhdl renameroo for output signals
  ap_cpu_data_master_requests_sdram_0_s1 <= internal_ap_cpu_data_master_requests_sdram_0_s1;
  --vhdl renameroo for output signals
  ap_cpu_instruction_master_granted_sdram_0_s1 <= internal_ap_cpu_instruction_master_granted_sdram_0_s1;
  --vhdl renameroo for output signals
  ap_cpu_instruction_master_qualified_request_sdram_0_s1 <= internal_ap_cpu_instruction_master_qualified_request_sdram_0_s1;
  --vhdl renameroo for output signals
  ap_cpu_instruction_master_requests_sdram_0_s1 <= internal_ap_cpu_instruction_master_requests_sdram_0_s1;
  --vhdl renameroo for output signals
  sdram_0_s1_waitrequest_from_sa <= internal_sdram_0_s1_waitrequest_from_sa;
--synthesis translate_off
    --sdram_0/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --grant signals are active simultaneously, which is an e_process
    process (clk)
    VARIABLE write_line47 : line;
    begin
      if clk'event and clk = '1' then
        if (std_logic_vector'("000000000000000000000000000000") & (((std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(internal_ap_cpu_data_master_granted_sdram_0_s1))) + (std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(internal_ap_cpu_instruction_master_granted_sdram_0_s1))))))>std_logic_vector'("00000000000000000000000000000001") then 
          write(write_line47, now);
          write(write_line47, string'(": "));
          write(write_line47, string'("> 1 of grant signals are active simultaneously"));
          write(output, write_line47.all);
          deallocate (write_line47);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --saved_grant signals are active simultaneously, which is an e_process
    process (clk)
    VARIABLE write_line48 : line;
    begin
      if clk'event and clk = '1' then
        if (std_logic_vector'("000000000000000000000000000000") & (((std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(ap_cpu_data_master_saved_grant_sdram_0_s1))) + (std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(ap_cpu_instruction_master_saved_grant_sdram_0_s1))))))>std_logic_vector'("00000000000000000000000000000001") then 
          write(write_line48, now);
          write(write_line48, string'(": "));
          write(write_line48, string'("> 1 of saved_grant signals are active simultaneously"));
          write(output, write_line48.all);
          deallocate (write_line48);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity status_led_pio_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal clock_crossing_0_m1_address_to_slave : IN STD_LOGIC_VECTOR (6 DOWNTO 0);
                 signal clock_crossing_0_m1_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal clock_crossing_0_m1_latency_counter : IN STD_LOGIC;
                 signal clock_crossing_0_m1_nativeaddress : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
                 signal clock_crossing_0_m1_read : IN STD_LOGIC;
                 signal clock_crossing_0_m1_write : IN STD_LOGIC;
                 signal clock_crossing_0_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;
                 signal status_led_pio_s1_readdata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);

              -- outputs:
                 signal clock_crossing_0_m1_granted_status_led_pio_s1 : OUT STD_LOGIC;
                 signal clock_crossing_0_m1_qualified_request_status_led_pio_s1 : OUT STD_LOGIC;
                 signal clock_crossing_0_m1_read_data_valid_status_led_pio_s1 : OUT STD_LOGIC;
                 signal clock_crossing_0_m1_requests_status_led_pio_s1 : OUT STD_LOGIC;
                 signal d1_status_led_pio_s1_end_xfer : OUT STD_LOGIC;
                 signal status_led_pio_s1_address : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal status_led_pio_s1_chipselect : OUT STD_LOGIC;
                 signal status_led_pio_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal status_led_pio_s1_reset_n : OUT STD_LOGIC;
                 signal status_led_pio_s1_write_n : OUT STD_LOGIC;
                 signal status_led_pio_s1_writedata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
              );
end entity status_led_pio_s1_arbitrator;


architecture europa of status_led_pio_s1_arbitrator is
                signal clock_crossing_0_m1_arbiterlock :  STD_LOGIC;
                signal clock_crossing_0_m1_arbiterlock2 :  STD_LOGIC;
                signal clock_crossing_0_m1_continuerequest :  STD_LOGIC;
                signal clock_crossing_0_m1_saved_grant_status_led_pio_s1 :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_status_led_pio_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_clock_crossing_0_m1_granted_status_led_pio_s1 :  STD_LOGIC;
                signal internal_clock_crossing_0_m1_qualified_request_status_led_pio_s1 :  STD_LOGIC;
                signal internal_clock_crossing_0_m1_requests_status_led_pio_s1 :  STD_LOGIC;
                signal status_led_pio_s1_allgrants :  STD_LOGIC;
                signal status_led_pio_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal status_led_pio_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal status_led_pio_s1_any_continuerequest :  STD_LOGIC;
                signal status_led_pio_s1_arb_counter_enable :  STD_LOGIC;
                signal status_led_pio_s1_arb_share_counter :  STD_LOGIC;
                signal status_led_pio_s1_arb_share_counter_next_value :  STD_LOGIC;
                signal status_led_pio_s1_arb_share_set_values :  STD_LOGIC;
                signal status_led_pio_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal status_led_pio_s1_begins_xfer :  STD_LOGIC;
                signal status_led_pio_s1_end_xfer :  STD_LOGIC;
                signal status_led_pio_s1_firsttransfer :  STD_LOGIC;
                signal status_led_pio_s1_grant_vector :  STD_LOGIC;
                signal status_led_pio_s1_in_a_read_cycle :  STD_LOGIC;
                signal status_led_pio_s1_in_a_write_cycle :  STD_LOGIC;
                signal status_led_pio_s1_master_qreq_vector :  STD_LOGIC;
                signal status_led_pio_s1_non_bursting_master_requests :  STD_LOGIC;
                signal status_led_pio_s1_pretend_byte_enable :  STD_LOGIC;
                signal status_led_pio_s1_reg_firsttransfer :  STD_LOGIC;
                signal status_led_pio_s1_slavearbiterlockenable :  STD_LOGIC;
                signal status_led_pio_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal status_led_pio_s1_unreg_firsttransfer :  STD_LOGIC;
                signal status_led_pio_s1_waits_for_read :  STD_LOGIC;
                signal status_led_pio_s1_waits_for_write :  STD_LOGIC;
                signal wait_for_status_led_pio_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT status_led_pio_s1_end_xfer;
    end if;

  end process;

  status_led_pio_s1_begins_xfer <= NOT d1_reasons_to_wait AND (internal_clock_crossing_0_m1_qualified_request_status_led_pio_s1);
  --assign status_led_pio_s1_readdata_from_sa = status_led_pio_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  status_led_pio_s1_readdata_from_sa <= status_led_pio_s1_readdata;
  internal_clock_crossing_0_m1_requests_status_led_pio_s1 <= to_std_logic(((Std_Logic_Vector'(clock_crossing_0_m1_address_to_slave(6 DOWNTO 5) & std_logic_vector'("00000")) = std_logic_vector'("0100000")))) AND ((clock_crossing_0_m1_read OR clock_crossing_0_m1_write));
  --status_led_pio_s1_arb_share_counter set values, which is an e_mux
  status_led_pio_s1_arb_share_set_values <= std_logic'('1');
  --status_led_pio_s1_non_bursting_master_requests mux, which is an e_mux
  status_led_pio_s1_non_bursting_master_requests <= internal_clock_crossing_0_m1_requests_status_led_pio_s1;
  --status_led_pio_s1_any_bursting_master_saved_grant mux, which is an e_mux
  status_led_pio_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --status_led_pio_s1_arb_share_counter_next_value assignment, which is an e_assign
  status_led_pio_s1_arb_share_counter_next_value <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(status_led_pio_s1_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(status_led_pio_s1_arb_share_set_values))) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(status_led_pio_s1_arb_share_counter) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(status_led_pio_s1_arb_share_counter))) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))));
  --status_led_pio_s1_allgrants all slave grants, which is an e_mux
  status_led_pio_s1_allgrants <= status_led_pio_s1_grant_vector;
  --status_led_pio_s1_end_xfer assignment, which is an e_assign
  status_led_pio_s1_end_xfer <= NOT ((status_led_pio_s1_waits_for_read OR status_led_pio_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_status_led_pio_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_status_led_pio_s1 <= status_led_pio_s1_end_xfer AND (((NOT status_led_pio_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --status_led_pio_s1_arb_share_counter arbitration counter enable, which is an e_assign
  status_led_pio_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_status_led_pio_s1 AND status_led_pio_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_status_led_pio_s1 AND NOT status_led_pio_s1_non_bursting_master_requests));
  --status_led_pio_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      status_led_pio_s1_arb_share_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(status_led_pio_s1_arb_counter_enable) = '1' then 
        status_led_pio_s1_arb_share_counter <= status_led_pio_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --status_led_pio_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      status_led_pio_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((status_led_pio_s1_master_qreq_vector AND end_xfer_arb_share_counter_term_status_led_pio_s1)) OR ((end_xfer_arb_share_counter_term_status_led_pio_s1 AND NOT status_led_pio_s1_non_bursting_master_requests)))) = '1' then 
        status_led_pio_s1_slavearbiterlockenable <= status_led_pio_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --clock_crossing_0/m1 status_led_pio/s1 arbiterlock, which is an e_assign
  clock_crossing_0_m1_arbiterlock <= status_led_pio_s1_slavearbiterlockenable AND clock_crossing_0_m1_continuerequest;
  --status_led_pio_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  status_led_pio_s1_slavearbiterlockenable2 <= status_led_pio_s1_arb_share_counter_next_value;
  --clock_crossing_0/m1 status_led_pio/s1 arbiterlock2, which is an e_assign
  clock_crossing_0_m1_arbiterlock2 <= status_led_pio_s1_slavearbiterlockenable2 AND clock_crossing_0_m1_continuerequest;
  --status_led_pio_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  status_led_pio_s1_any_continuerequest <= std_logic'('1');
  --clock_crossing_0_m1_continuerequest continued request, which is an e_assign
  clock_crossing_0_m1_continuerequest <= std_logic'('1');
  internal_clock_crossing_0_m1_qualified_request_status_led_pio_s1 <= internal_clock_crossing_0_m1_requests_status_led_pio_s1 AND NOT ((clock_crossing_0_m1_read AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(clock_crossing_0_m1_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))))));
  --local readdatavalid clock_crossing_0_m1_read_data_valid_status_led_pio_s1, which is an e_mux
  clock_crossing_0_m1_read_data_valid_status_led_pio_s1 <= (internal_clock_crossing_0_m1_granted_status_led_pio_s1 AND clock_crossing_0_m1_read) AND NOT status_led_pio_s1_waits_for_read;
  --status_led_pio_s1_writedata mux, which is an e_mux
  status_led_pio_s1_writedata <= clock_crossing_0_m1_writedata (7 DOWNTO 0);
  --master is always granted when requested
  internal_clock_crossing_0_m1_granted_status_led_pio_s1 <= internal_clock_crossing_0_m1_qualified_request_status_led_pio_s1;
  --clock_crossing_0/m1 saved-grant status_led_pio/s1, which is an e_assign
  clock_crossing_0_m1_saved_grant_status_led_pio_s1 <= internal_clock_crossing_0_m1_requests_status_led_pio_s1;
  --allow new arb cycle for status_led_pio/s1, which is an e_assign
  status_led_pio_s1_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  status_led_pio_s1_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  status_led_pio_s1_master_qreq_vector <= std_logic'('1');
  --status_led_pio_s1_reset_n assignment, which is an e_assign
  status_led_pio_s1_reset_n <= reset_n;
  status_led_pio_s1_chipselect <= internal_clock_crossing_0_m1_granted_status_led_pio_s1;
  --status_led_pio_s1_firsttransfer first transaction, which is an e_assign
  status_led_pio_s1_firsttransfer <= A_WE_StdLogic((std_logic'(status_led_pio_s1_begins_xfer) = '1'), status_led_pio_s1_unreg_firsttransfer, status_led_pio_s1_reg_firsttransfer);
  --status_led_pio_s1_unreg_firsttransfer first transaction, which is an e_assign
  status_led_pio_s1_unreg_firsttransfer <= NOT ((status_led_pio_s1_slavearbiterlockenable AND status_led_pio_s1_any_continuerequest));
  --status_led_pio_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      status_led_pio_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(status_led_pio_s1_begins_xfer) = '1' then 
        status_led_pio_s1_reg_firsttransfer <= status_led_pio_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --status_led_pio_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  status_led_pio_s1_beginbursttransfer_internal <= status_led_pio_s1_begins_xfer;
  --~status_led_pio_s1_write_n assignment, which is an e_mux
  status_led_pio_s1_write_n <= NOT ((((internal_clock_crossing_0_m1_granted_status_led_pio_s1 AND clock_crossing_0_m1_write)) AND status_led_pio_s1_pretend_byte_enable));
  --status_led_pio_s1_address mux, which is an e_mux
  status_led_pio_s1_address <= clock_crossing_0_m1_nativeaddress (2 DOWNTO 0);
  --d1_status_led_pio_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_status_led_pio_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_status_led_pio_s1_end_xfer <= status_led_pio_s1_end_xfer;
    end if;

  end process;

  --status_led_pio_s1_waits_for_read in a cycle, which is an e_mux
  status_led_pio_s1_waits_for_read <= status_led_pio_s1_in_a_read_cycle AND status_led_pio_s1_begins_xfer;
  --status_led_pio_s1_in_a_read_cycle assignment, which is an e_assign
  status_led_pio_s1_in_a_read_cycle <= internal_clock_crossing_0_m1_granted_status_led_pio_s1 AND clock_crossing_0_m1_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= status_led_pio_s1_in_a_read_cycle;
  --status_led_pio_s1_waits_for_write in a cycle, which is an e_mux
  status_led_pio_s1_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(status_led_pio_s1_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --status_led_pio_s1_in_a_write_cycle assignment, which is an e_assign
  status_led_pio_s1_in_a_write_cycle <= internal_clock_crossing_0_m1_granted_status_led_pio_s1 AND clock_crossing_0_m1_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= status_led_pio_s1_in_a_write_cycle;
  wait_for_status_led_pio_s1_counter <= std_logic'('0');
  --status_led_pio_s1_pretend_byte_enable byte enable port mux, which is an e_mux
  status_led_pio_s1_pretend_byte_enable <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((internal_clock_crossing_0_m1_granted_status_led_pio_s1)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (clock_crossing_0_m1_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))));
  --vhdl renameroo for output signals
  clock_crossing_0_m1_granted_status_led_pio_s1 <= internal_clock_crossing_0_m1_granted_status_led_pio_s1;
  --vhdl renameroo for output signals
  clock_crossing_0_m1_qualified_request_status_led_pio_s1 <= internal_clock_crossing_0_m1_qualified_request_status_led_pio_s1;
  --vhdl renameroo for output signals
  clock_crossing_0_m1_requests_status_led_pio_s1 <= internal_clock_crossing_0_m1_requests_status_led_pio_s1;
--synthesis translate_off
    --status_led_pio/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity sync_irq_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal clock_crossing_1_m1_address_to_slave : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal clock_crossing_1_m1_latency_counter : IN STD_LOGIC;
                 signal clock_crossing_1_m1_nativeaddress : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
                 signal clock_crossing_1_m1_read : IN STD_LOGIC;
                 signal clock_crossing_1_m1_write : IN STD_LOGIC;
                 signal clock_crossing_1_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;
                 signal sync_irq_s1_irq : IN STD_LOGIC;
                 signal sync_irq_s1_readdata : IN STD_LOGIC;

              -- outputs:
                 signal clock_crossing_1_m1_granted_sync_irq_s1 : OUT STD_LOGIC;
                 signal clock_crossing_1_m1_qualified_request_sync_irq_s1 : OUT STD_LOGIC;
                 signal clock_crossing_1_m1_read_data_valid_sync_irq_s1 : OUT STD_LOGIC;
                 signal clock_crossing_1_m1_requests_sync_irq_s1 : OUT STD_LOGIC;
                 signal d1_sync_irq_s1_end_xfer : OUT STD_LOGIC;
                 signal sync_irq_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal sync_irq_s1_chipselect : OUT STD_LOGIC;
                 signal sync_irq_s1_irq_from_sa : OUT STD_LOGIC;
                 signal sync_irq_s1_readdata_from_sa : OUT STD_LOGIC;
                 signal sync_irq_s1_reset_n : OUT STD_LOGIC;
                 signal sync_irq_s1_write_n : OUT STD_LOGIC;
                 signal sync_irq_s1_writedata : OUT STD_LOGIC
              );
end entity sync_irq_s1_arbitrator;


architecture europa of sync_irq_s1_arbitrator is
                signal clock_crossing_1_m1_arbiterlock :  STD_LOGIC;
                signal clock_crossing_1_m1_arbiterlock2 :  STD_LOGIC;
                signal clock_crossing_1_m1_continuerequest :  STD_LOGIC;
                signal clock_crossing_1_m1_saved_grant_sync_irq_s1 :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_sync_irq_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_clock_crossing_1_m1_granted_sync_irq_s1 :  STD_LOGIC;
                signal internal_clock_crossing_1_m1_qualified_request_sync_irq_s1 :  STD_LOGIC;
                signal internal_clock_crossing_1_m1_requests_sync_irq_s1 :  STD_LOGIC;
                signal sync_irq_s1_allgrants :  STD_LOGIC;
                signal sync_irq_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal sync_irq_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal sync_irq_s1_any_continuerequest :  STD_LOGIC;
                signal sync_irq_s1_arb_counter_enable :  STD_LOGIC;
                signal sync_irq_s1_arb_share_counter :  STD_LOGIC;
                signal sync_irq_s1_arb_share_counter_next_value :  STD_LOGIC;
                signal sync_irq_s1_arb_share_set_values :  STD_LOGIC;
                signal sync_irq_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal sync_irq_s1_begins_xfer :  STD_LOGIC;
                signal sync_irq_s1_end_xfer :  STD_LOGIC;
                signal sync_irq_s1_firsttransfer :  STD_LOGIC;
                signal sync_irq_s1_grant_vector :  STD_LOGIC;
                signal sync_irq_s1_in_a_read_cycle :  STD_LOGIC;
                signal sync_irq_s1_in_a_write_cycle :  STD_LOGIC;
                signal sync_irq_s1_master_qreq_vector :  STD_LOGIC;
                signal sync_irq_s1_non_bursting_master_requests :  STD_LOGIC;
                signal sync_irq_s1_reg_firsttransfer :  STD_LOGIC;
                signal sync_irq_s1_slavearbiterlockenable :  STD_LOGIC;
                signal sync_irq_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal sync_irq_s1_unreg_firsttransfer :  STD_LOGIC;
                signal sync_irq_s1_waits_for_read :  STD_LOGIC;
                signal sync_irq_s1_waits_for_write :  STD_LOGIC;
                signal wait_for_sync_irq_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT sync_irq_s1_end_xfer;
    end if;

  end process;

  sync_irq_s1_begins_xfer <= NOT d1_reasons_to_wait AND (internal_clock_crossing_1_m1_qualified_request_sync_irq_s1);
  --assign sync_irq_s1_readdata_from_sa = sync_irq_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  sync_irq_s1_readdata_from_sa <= sync_irq_s1_readdata;
  internal_clock_crossing_1_m1_requests_sync_irq_s1 <= to_std_logic(((Std_Logic_Vector'(clock_crossing_1_m1_address_to_slave(7 DOWNTO 4) & std_logic_vector'("0000")) = std_logic_vector'("11000000")))) AND ((clock_crossing_1_m1_read OR clock_crossing_1_m1_write));
  --sync_irq_s1_arb_share_counter set values, which is an e_mux
  sync_irq_s1_arb_share_set_values <= std_logic'('1');
  --sync_irq_s1_non_bursting_master_requests mux, which is an e_mux
  sync_irq_s1_non_bursting_master_requests <= internal_clock_crossing_1_m1_requests_sync_irq_s1;
  --sync_irq_s1_any_bursting_master_saved_grant mux, which is an e_mux
  sync_irq_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --sync_irq_s1_arb_share_counter_next_value assignment, which is an e_assign
  sync_irq_s1_arb_share_counter_next_value <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(sync_irq_s1_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(sync_irq_s1_arb_share_set_values))) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(sync_irq_s1_arb_share_counter) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(sync_irq_s1_arb_share_counter))) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))));
  --sync_irq_s1_allgrants all slave grants, which is an e_mux
  sync_irq_s1_allgrants <= sync_irq_s1_grant_vector;
  --sync_irq_s1_end_xfer assignment, which is an e_assign
  sync_irq_s1_end_xfer <= NOT ((sync_irq_s1_waits_for_read OR sync_irq_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_sync_irq_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_sync_irq_s1 <= sync_irq_s1_end_xfer AND (((NOT sync_irq_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --sync_irq_s1_arb_share_counter arbitration counter enable, which is an e_assign
  sync_irq_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_sync_irq_s1 AND sync_irq_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_sync_irq_s1 AND NOT sync_irq_s1_non_bursting_master_requests));
  --sync_irq_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sync_irq_s1_arb_share_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(sync_irq_s1_arb_counter_enable) = '1' then 
        sync_irq_s1_arb_share_counter <= sync_irq_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --sync_irq_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sync_irq_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((sync_irq_s1_master_qreq_vector AND end_xfer_arb_share_counter_term_sync_irq_s1)) OR ((end_xfer_arb_share_counter_term_sync_irq_s1 AND NOT sync_irq_s1_non_bursting_master_requests)))) = '1' then 
        sync_irq_s1_slavearbiterlockenable <= sync_irq_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --clock_crossing_1/m1 sync_irq/s1 arbiterlock, which is an e_assign
  clock_crossing_1_m1_arbiterlock <= sync_irq_s1_slavearbiterlockenable AND clock_crossing_1_m1_continuerequest;
  --sync_irq_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  sync_irq_s1_slavearbiterlockenable2 <= sync_irq_s1_arb_share_counter_next_value;
  --clock_crossing_1/m1 sync_irq/s1 arbiterlock2, which is an e_assign
  clock_crossing_1_m1_arbiterlock2 <= sync_irq_s1_slavearbiterlockenable2 AND clock_crossing_1_m1_continuerequest;
  --sync_irq_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  sync_irq_s1_any_continuerequest <= std_logic'('1');
  --clock_crossing_1_m1_continuerequest continued request, which is an e_assign
  clock_crossing_1_m1_continuerequest <= std_logic'('1');
  internal_clock_crossing_1_m1_qualified_request_sync_irq_s1 <= internal_clock_crossing_1_m1_requests_sync_irq_s1 AND NOT ((clock_crossing_1_m1_read AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(clock_crossing_1_m1_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))))));
  --local readdatavalid clock_crossing_1_m1_read_data_valid_sync_irq_s1, which is an e_mux
  clock_crossing_1_m1_read_data_valid_sync_irq_s1 <= (internal_clock_crossing_1_m1_granted_sync_irq_s1 AND clock_crossing_1_m1_read) AND NOT sync_irq_s1_waits_for_read;
  --sync_irq_s1_writedata mux, which is an e_mux
  sync_irq_s1_writedata <= clock_crossing_1_m1_writedata(0);
  --master is always granted when requested
  internal_clock_crossing_1_m1_granted_sync_irq_s1 <= internal_clock_crossing_1_m1_qualified_request_sync_irq_s1;
  --clock_crossing_1/m1 saved-grant sync_irq/s1, which is an e_assign
  clock_crossing_1_m1_saved_grant_sync_irq_s1 <= internal_clock_crossing_1_m1_requests_sync_irq_s1;
  --allow new arb cycle for sync_irq/s1, which is an e_assign
  sync_irq_s1_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  sync_irq_s1_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  sync_irq_s1_master_qreq_vector <= std_logic'('1');
  --sync_irq_s1_reset_n assignment, which is an e_assign
  sync_irq_s1_reset_n <= reset_n;
  sync_irq_s1_chipselect <= internal_clock_crossing_1_m1_granted_sync_irq_s1;
  --sync_irq_s1_firsttransfer first transaction, which is an e_assign
  sync_irq_s1_firsttransfer <= A_WE_StdLogic((std_logic'(sync_irq_s1_begins_xfer) = '1'), sync_irq_s1_unreg_firsttransfer, sync_irq_s1_reg_firsttransfer);
  --sync_irq_s1_unreg_firsttransfer first transaction, which is an e_assign
  sync_irq_s1_unreg_firsttransfer <= NOT ((sync_irq_s1_slavearbiterlockenable AND sync_irq_s1_any_continuerequest));
  --sync_irq_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sync_irq_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(sync_irq_s1_begins_xfer) = '1' then 
        sync_irq_s1_reg_firsttransfer <= sync_irq_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --sync_irq_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  sync_irq_s1_beginbursttransfer_internal <= sync_irq_s1_begins_xfer;
  --~sync_irq_s1_write_n assignment, which is an e_mux
  sync_irq_s1_write_n <= NOT ((internal_clock_crossing_1_m1_granted_sync_irq_s1 AND clock_crossing_1_m1_write));
  --sync_irq_s1_address mux, which is an e_mux
  sync_irq_s1_address <= clock_crossing_1_m1_nativeaddress (1 DOWNTO 0);
  --d1_sync_irq_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_sync_irq_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_sync_irq_s1_end_xfer <= sync_irq_s1_end_xfer;
    end if;

  end process;

  --sync_irq_s1_waits_for_read in a cycle, which is an e_mux
  sync_irq_s1_waits_for_read <= sync_irq_s1_in_a_read_cycle AND sync_irq_s1_begins_xfer;
  --sync_irq_s1_in_a_read_cycle assignment, which is an e_assign
  sync_irq_s1_in_a_read_cycle <= internal_clock_crossing_1_m1_granted_sync_irq_s1 AND clock_crossing_1_m1_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= sync_irq_s1_in_a_read_cycle;
  --sync_irq_s1_waits_for_write in a cycle, which is an e_mux
  sync_irq_s1_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(sync_irq_s1_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --sync_irq_s1_in_a_write_cycle assignment, which is an e_assign
  sync_irq_s1_in_a_write_cycle <= internal_clock_crossing_1_m1_granted_sync_irq_s1 AND clock_crossing_1_m1_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= sync_irq_s1_in_a_write_cycle;
  wait_for_sync_irq_s1_counter <= std_logic'('0');
  --assign sync_irq_s1_irq_from_sa = sync_irq_s1_irq so that symbol knows where to group signals which may go to master only, which is an e_assign
  sync_irq_s1_irq_from_sa <= sync_irq_s1_irq;
  --vhdl renameroo for output signals
  clock_crossing_1_m1_granted_sync_irq_s1 <= internal_clock_crossing_1_m1_granted_sync_irq_s1;
  --vhdl renameroo for output signals
  clock_crossing_1_m1_qualified_request_sync_irq_s1 <= internal_clock_crossing_1_m1_qualified_request_sync_irq_s1;
  --vhdl renameroo for output signals
  clock_crossing_1_m1_requests_sync_irq_s1 <= internal_clock_crossing_1_m1_requests_sync_irq_s1;
--synthesis translate_off
    --sync_irq/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity sysid_control_slave_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal clock_crossing_0_m1_address_to_slave : IN STD_LOGIC_VECTOR (6 DOWNTO 0);
                 signal clock_crossing_0_m1_latency_counter : IN STD_LOGIC;
                 signal clock_crossing_0_m1_nativeaddress : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
                 signal clock_crossing_0_m1_read : IN STD_LOGIC;
                 signal clock_crossing_0_m1_write : IN STD_LOGIC;
                 signal clock_crossing_1_m1_address_to_slave : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal clock_crossing_1_m1_latency_counter : IN STD_LOGIC;
                 signal clock_crossing_1_m1_nativeaddress : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
                 signal clock_crossing_1_m1_read : IN STD_LOGIC;
                 signal clock_crossing_1_m1_write : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sysid_control_slave_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

              -- outputs:
                 signal clock_crossing_0_m1_granted_sysid_control_slave : OUT STD_LOGIC;
                 signal clock_crossing_0_m1_qualified_request_sysid_control_slave : OUT STD_LOGIC;
                 signal clock_crossing_0_m1_read_data_valid_sysid_control_slave : OUT STD_LOGIC;
                 signal clock_crossing_0_m1_requests_sysid_control_slave : OUT STD_LOGIC;
                 signal clock_crossing_1_m1_granted_sysid_control_slave : OUT STD_LOGIC;
                 signal clock_crossing_1_m1_qualified_request_sysid_control_slave : OUT STD_LOGIC;
                 signal clock_crossing_1_m1_read_data_valid_sysid_control_slave : OUT STD_LOGIC;
                 signal clock_crossing_1_m1_requests_sysid_control_slave : OUT STD_LOGIC;
                 signal d1_sysid_control_slave_end_xfer : OUT STD_LOGIC;
                 signal sysid_control_slave_address : OUT STD_LOGIC;
                 signal sysid_control_slave_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
              );
end entity sysid_control_slave_arbitrator;


architecture europa of sysid_control_slave_arbitrator is
                signal clock_crossing_0_m1_arbiterlock :  STD_LOGIC;
                signal clock_crossing_0_m1_arbiterlock2 :  STD_LOGIC;
                signal clock_crossing_0_m1_continuerequest :  STD_LOGIC;
                signal clock_crossing_0_m1_saved_grant_sysid_control_slave :  STD_LOGIC;
                signal clock_crossing_1_m1_arbiterlock :  STD_LOGIC;
                signal clock_crossing_1_m1_arbiterlock2 :  STD_LOGIC;
                signal clock_crossing_1_m1_continuerequest :  STD_LOGIC;
                signal clock_crossing_1_m1_saved_grant_sysid_control_slave :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_sysid_control_slave :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_clock_crossing_0_m1_granted_sysid_control_slave :  STD_LOGIC;
                signal internal_clock_crossing_0_m1_qualified_request_sysid_control_slave :  STD_LOGIC;
                signal internal_clock_crossing_0_m1_requests_sysid_control_slave :  STD_LOGIC;
                signal internal_clock_crossing_1_m1_granted_sysid_control_slave :  STD_LOGIC;
                signal internal_clock_crossing_1_m1_qualified_request_sysid_control_slave :  STD_LOGIC;
                signal internal_clock_crossing_1_m1_requests_sysid_control_slave :  STD_LOGIC;
                signal last_cycle_clock_crossing_0_m1_granted_slave_sysid_control_slave :  STD_LOGIC;
                signal last_cycle_clock_crossing_1_m1_granted_slave_sysid_control_slave :  STD_LOGIC;
                signal sysid_control_slave_allgrants :  STD_LOGIC;
                signal sysid_control_slave_allow_new_arb_cycle :  STD_LOGIC;
                signal sysid_control_slave_any_bursting_master_saved_grant :  STD_LOGIC;
                signal sysid_control_slave_any_continuerequest :  STD_LOGIC;
                signal sysid_control_slave_arb_addend :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal sysid_control_slave_arb_counter_enable :  STD_LOGIC;
                signal sysid_control_slave_arb_share_counter :  STD_LOGIC;
                signal sysid_control_slave_arb_share_counter_next_value :  STD_LOGIC;
                signal sysid_control_slave_arb_share_set_values :  STD_LOGIC;
                signal sysid_control_slave_arb_winner :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal sysid_control_slave_arbitration_holdoff_internal :  STD_LOGIC;
                signal sysid_control_slave_beginbursttransfer_internal :  STD_LOGIC;
                signal sysid_control_slave_begins_xfer :  STD_LOGIC;
                signal sysid_control_slave_chosen_master_double_vector :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal sysid_control_slave_chosen_master_rot_left :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal sysid_control_slave_end_xfer :  STD_LOGIC;
                signal sysid_control_slave_firsttransfer :  STD_LOGIC;
                signal sysid_control_slave_grant_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal sysid_control_slave_in_a_read_cycle :  STD_LOGIC;
                signal sysid_control_slave_in_a_write_cycle :  STD_LOGIC;
                signal sysid_control_slave_master_qreq_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal sysid_control_slave_non_bursting_master_requests :  STD_LOGIC;
                signal sysid_control_slave_reg_firsttransfer :  STD_LOGIC;
                signal sysid_control_slave_saved_chosen_master_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal sysid_control_slave_slavearbiterlockenable :  STD_LOGIC;
                signal sysid_control_slave_slavearbiterlockenable2 :  STD_LOGIC;
                signal sysid_control_slave_unreg_firsttransfer :  STD_LOGIC;
                signal sysid_control_slave_waits_for_read :  STD_LOGIC;
                signal sysid_control_slave_waits_for_write :  STD_LOGIC;
                signal wait_for_sysid_control_slave_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT sysid_control_slave_end_xfer;
    end if;

  end process;

  sysid_control_slave_begins_xfer <= NOT d1_reasons_to_wait AND ((internal_clock_crossing_0_m1_qualified_request_sysid_control_slave OR internal_clock_crossing_1_m1_qualified_request_sysid_control_slave));
  --assign sysid_control_slave_readdata_from_sa = sysid_control_slave_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  sysid_control_slave_readdata_from_sa <= sysid_control_slave_readdata;
  internal_clock_crossing_0_m1_requests_sysid_control_slave <= ((to_std_logic(((Std_Logic_Vector'(clock_crossing_0_m1_address_to_slave(6 DOWNTO 3) & std_logic_vector'("000")) = std_logic_vector'("1100000")))) AND ((clock_crossing_0_m1_read OR clock_crossing_0_m1_write)))) AND clock_crossing_0_m1_read;
  --sysid_control_slave_arb_share_counter set values, which is an e_mux
  sysid_control_slave_arb_share_set_values <= std_logic'('1');
  --sysid_control_slave_non_bursting_master_requests mux, which is an e_mux
  sysid_control_slave_non_bursting_master_requests <= ((internal_clock_crossing_0_m1_requests_sysid_control_slave OR internal_clock_crossing_1_m1_requests_sysid_control_slave) OR internal_clock_crossing_0_m1_requests_sysid_control_slave) OR internal_clock_crossing_1_m1_requests_sysid_control_slave;
  --sysid_control_slave_any_bursting_master_saved_grant mux, which is an e_mux
  sysid_control_slave_any_bursting_master_saved_grant <= std_logic'('0');
  --sysid_control_slave_arb_share_counter_next_value assignment, which is an e_assign
  sysid_control_slave_arb_share_counter_next_value <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(sysid_control_slave_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(sysid_control_slave_arb_share_set_values))) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(sysid_control_slave_arb_share_counter) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(sysid_control_slave_arb_share_counter))) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))));
  --sysid_control_slave_allgrants all slave grants, which is an e_mux
  sysid_control_slave_allgrants <= (((or_reduce(sysid_control_slave_grant_vector)) OR (or_reduce(sysid_control_slave_grant_vector))) OR (or_reduce(sysid_control_slave_grant_vector))) OR (or_reduce(sysid_control_slave_grant_vector));
  --sysid_control_slave_end_xfer assignment, which is an e_assign
  sysid_control_slave_end_xfer <= NOT ((sysid_control_slave_waits_for_read OR sysid_control_slave_waits_for_write));
  --end_xfer_arb_share_counter_term_sysid_control_slave arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_sysid_control_slave <= sysid_control_slave_end_xfer AND (((NOT sysid_control_slave_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --sysid_control_slave_arb_share_counter arbitration counter enable, which is an e_assign
  sysid_control_slave_arb_counter_enable <= ((end_xfer_arb_share_counter_term_sysid_control_slave AND sysid_control_slave_allgrants)) OR ((end_xfer_arb_share_counter_term_sysid_control_slave AND NOT sysid_control_slave_non_bursting_master_requests));
  --sysid_control_slave_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sysid_control_slave_arb_share_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(sysid_control_slave_arb_counter_enable) = '1' then 
        sysid_control_slave_arb_share_counter <= sysid_control_slave_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --sysid_control_slave_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sysid_control_slave_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((or_reduce(sysid_control_slave_master_qreq_vector) AND end_xfer_arb_share_counter_term_sysid_control_slave)) OR ((end_xfer_arb_share_counter_term_sysid_control_slave AND NOT sysid_control_slave_non_bursting_master_requests)))) = '1' then 
        sysid_control_slave_slavearbiterlockenable <= sysid_control_slave_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --clock_crossing_0/m1 sysid/control_slave arbiterlock, which is an e_assign
  clock_crossing_0_m1_arbiterlock <= sysid_control_slave_slavearbiterlockenable AND clock_crossing_0_m1_continuerequest;
  --sysid_control_slave_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  sysid_control_slave_slavearbiterlockenable2 <= sysid_control_slave_arb_share_counter_next_value;
  --clock_crossing_0/m1 sysid/control_slave arbiterlock2, which is an e_assign
  clock_crossing_0_m1_arbiterlock2 <= sysid_control_slave_slavearbiterlockenable2 AND clock_crossing_0_m1_continuerequest;
  --clock_crossing_1/m1 sysid/control_slave arbiterlock, which is an e_assign
  clock_crossing_1_m1_arbiterlock <= sysid_control_slave_slavearbiterlockenable AND clock_crossing_1_m1_continuerequest;
  --clock_crossing_1/m1 sysid/control_slave arbiterlock2, which is an e_assign
  clock_crossing_1_m1_arbiterlock2 <= sysid_control_slave_slavearbiterlockenable2 AND clock_crossing_1_m1_continuerequest;
  --clock_crossing_1/m1 granted sysid/control_slave last time, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      last_cycle_clock_crossing_1_m1_granted_slave_sysid_control_slave <= std_logic'('0');
    elsif clk'event and clk = '1' then
      last_cycle_clock_crossing_1_m1_granted_slave_sysid_control_slave <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(clock_crossing_1_m1_saved_grant_sysid_control_slave) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((sysid_control_slave_arbitration_holdoff_internal OR NOT internal_clock_crossing_1_m1_requests_sysid_control_slave))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_clock_crossing_1_m1_granted_slave_sysid_control_slave))))));
    end if;

  end process;

  --clock_crossing_1_m1_continuerequest continued request, which is an e_mux
  clock_crossing_1_m1_continuerequest <= last_cycle_clock_crossing_1_m1_granted_slave_sysid_control_slave AND internal_clock_crossing_1_m1_requests_sysid_control_slave;
  --sysid_control_slave_any_continuerequest at least one master continues requesting, which is an e_mux
  sysid_control_slave_any_continuerequest <= clock_crossing_1_m1_continuerequest OR clock_crossing_0_m1_continuerequest;
  internal_clock_crossing_0_m1_qualified_request_sysid_control_slave <= internal_clock_crossing_0_m1_requests_sysid_control_slave AND NOT ((((clock_crossing_0_m1_read AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(clock_crossing_0_m1_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000")))))) OR clock_crossing_1_m1_arbiterlock));
  --local readdatavalid clock_crossing_0_m1_read_data_valid_sysid_control_slave, which is an e_mux
  clock_crossing_0_m1_read_data_valid_sysid_control_slave <= (internal_clock_crossing_0_m1_granted_sysid_control_slave AND clock_crossing_0_m1_read) AND NOT sysid_control_slave_waits_for_read;
  internal_clock_crossing_1_m1_requests_sysid_control_slave <= ((to_std_logic(((Std_Logic_Vector'(clock_crossing_1_m1_address_to_slave(7 DOWNTO 3) & std_logic_vector'("000")) = std_logic_vector'("01100000")))) AND ((clock_crossing_1_m1_read OR clock_crossing_1_m1_write)))) AND clock_crossing_1_m1_read;
  --clock_crossing_0/m1 granted sysid/control_slave last time, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      last_cycle_clock_crossing_0_m1_granted_slave_sysid_control_slave <= std_logic'('0');
    elsif clk'event and clk = '1' then
      last_cycle_clock_crossing_0_m1_granted_slave_sysid_control_slave <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(clock_crossing_0_m1_saved_grant_sysid_control_slave) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((sysid_control_slave_arbitration_holdoff_internal OR NOT internal_clock_crossing_0_m1_requests_sysid_control_slave))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_clock_crossing_0_m1_granted_slave_sysid_control_slave))))));
    end if;

  end process;

  --clock_crossing_0_m1_continuerequest continued request, which is an e_mux
  clock_crossing_0_m1_continuerequest <= last_cycle_clock_crossing_0_m1_granted_slave_sysid_control_slave AND internal_clock_crossing_0_m1_requests_sysid_control_slave;
  internal_clock_crossing_1_m1_qualified_request_sysid_control_slave <= internal_clock_crossing_1_m1_requests_sysid_control_slave AND NOT ((((clock_crossing_1_m1_read AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(clock_crossing_1_m1_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000")))))) OR clock_crossing_0_m1_arbiterlock));
  --local readdatavalid clock_crossing_1_m1_read_data_valid_sysid_control_slave, which is an e_mux
  clock_crossing_1_m1_read_data_valid_sysid_control_slave <= (internal_clock_crossing_1_m1_granted_sysid_control_slave AND clock_crossing_1_m1_read) AND NOT sysid_control_slave_waits_for_read;
  --allow new arb cycle for sysid/control_slave, which is an e_assign
  sysid_control_slave_allow_new_arb_cycle <= NOT clock_crossing_0_m1_arbiterlock AND NOT clock_crossing_1_m1_arbiterlock;
  --clock_crossing_1/m1 assignment into master qualified-requests vector for sysid/control_slave, which is an e_assign
  sysid_control_slave_master_qreq_vector(0) <= internal_clock_crossing_1_m1_qualified_request_sysid_control_slave;
  --clock_crossing_1/m1 grant sysid/control_slave, which is an e_assign
  internal_clock_crossing_1_m1_granted_sysid_control_slave <= sysid_control_slave_grant_vector(0);
  --clock_crossing_1/m1 saved-grant sysid/control_slave, which is an e_assign
  clock_crossing_1_m1_saved_grant_sysid_control_slave <= sysid_control_slave_arb_winner(0) AND internal_clock_crossing_1_m1_requests_sysid_control_slave;
  --clock_crossing_0/m1 assignment into master qualified-requests vector for sysid/control_slave, which is an e_assign
  sysid_control_slave_master_qreq_vector(1) <= internal_clock_crossing_0_m1_qualified_request_sysid_control_slave;
  --clock_crossing_0/m1 grant sysid/control_slave, which is an e_assign
  internal_clock_crossing_0_m1_granted_sysid_control_slave <= sysid_control_slave_grant_vector(1);
  --clock_crossing_0/m1 saved-grant sysid/control_slave, which is an e_assign
  clock_crossing_0_m1_saved_grant_sysid_control_slave <= sysid_control_slave_arb_winner(1) AND internal_clock_crossing_0_m1_requests_sysid_control_slave;
  --sysid/control_slave chosen-master double-vector, which is an e_assign
  sysid_control_slave_chosen_master_double_vector <= A_EXT (((std_logic_vector'("0") & ((sysid_control_slave_master_qreq_vector & sysid_control_slave_master_qreq_vector))) AND (((std_logic_vector'("0") & (Std_Logic_Vector'(NOT sysid_control_slave_master_qreq_vector & NOT sysid_control_slave_master_qreq_vector))) + (std_logic_vector'("000") & (sysid_control_slave_arb_addend))))), 4);
  --stable onehot encoding of arb winner
  sysid_control_slave_arb_winner <= A_WE_StdLogicVector((std_logic'(((sysid_control_slave_allow_new_arb_cycle AND or_reduce(sysid_control_slave_grant_vector)))) = '1'), sysid_control_slave_grant_vector, sysid_control_slave_saved_chosen_master_vector);
  --saved sysid_control_slave_grant_vector, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sysid_control_slave_saved_chosen_master_vector <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      if std_logic'(sysid_control_slave_allow_new_arb_cycle) = '1' then 
        sysid_control_slave_saved_chosen_master_vector <= A_WE_StdLogicVector((std_logic'(or_reduce(sysid_control_slave_grant_vector)) = '1'), sysid_control_slave_grant_vector, sysid_control_slave_saved_chosen_master_vector);
      end if;
    end if;

  end process;

  --onehot encoding of chosen master
  sysid_control_slave_grant_vector <= Std_Logic_Vector'(A_ToStdLogicVector(((sysid_control_slave_chosen_master_double_vector(1) OR sysid_control_slave_chosen_master_double_vector(3)))) & A_ToStdLogicVector(((sysid_control_slave_chosen_master_double_vector(0) OR sysid_control_slave_chosen_master_double_vector(2)))));
  --sysid/control_slave chosen master rotated left, which is an e_assign
  sysid_control_slave_chosen_master_rot_left <= A_EXT (A_WE_StdLogicVector((((A_SLL(sysid_control_slave_arb_winner,std_logic_vector'("00000000000000000000000000000001")))) /= std_logic_vector'("00")), (std_logic_vector'("000000000000000000000000000000") & ((A_SLL(sysid_control_slave_arb_winner,std_logic_vector'("00000000000000000000000000000001"))))), std_logic_vector'("00000000000000000000000000000001")), 2);
  --sysid/control_slave's addend for next-master-grant
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sysid_control_slave_arb_addend <= std_logic_vector'("01");
    elsif clk'event and clk = '1' then
      if std_logic'(or_reduce(sysid_control_slave_grant_vector)) = '1' then 
        sysid_control_slave_arb_addend <= A_WE_StdLogicVector((std_logic'(sysid_control_slave_end_xfer) = '1'), sysid_control_slave_chosen_master_rot_left, sysid_control_slave_grant_vector);
      end if;
    end if;

  end process;

  --sysid_control_slave_firsttransfer first transaction, which is an e_assign
  sysid_control_slave_firsttransfer <= A_WE_StdLogic((std_logic'(sysid_control_slave_begins_xfer) = '1'), sysid_control_slave_unreg_firsttransfer, sysid_control_slave_reg_firsttransfer);
  --sysid_control_slave_unreg_firsttransfer first transaction, which is an e_assign
  sysid_control_slave_unreg_firsttransfer <= NOT ((sysid_control_slave_slavearbiterlockenable AND sysid_control_slave_any_continuerequest));
  --sysid_control_slave_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sysid_control_slave_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(sysid_control_slave_begins_xfer) = '1' then 
        sysid_control_slave_reg_firsttransfer <= sysid_control_slave_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --sysid_control_slave_beginbursttransfer_internal begin burst transfer, which is an e_assign
  sysid_control_slave_beginbursttransfer_internal <= sysid_control_slave_begins_xfer;
  --sysid_control_slave_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  sysid_control_slave_arbitration_holdoff_internal <= sysid_control_slave_begins_xfer AND sysid_control_slave_firsttransfer;
  --sysid_control_slave_address mux, which is an e_mux
  sysid_control_slave_address <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((internal_clock_crossing_0_m1_granted_sysid_control_slave)) = '1'), (std_logic_vector'("0") & (clock_crossing_0_m1_nativeaddress)), clock_crossing_1_m1_nativeaddress));
  --d1_sysid_control_slave_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_sysid_control_slave_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_sysid_control_slave_end_xfer <= sysid_control_slave_end_xfer;
    end if;

  end process;

  --sysid_control_slave_waits_for_read in a cycle, which is an e_mux
  sysid_control_slave_waits_for_read <= sysid_control_slave_in_a_read_cycle AND sysid_control_slave_begins_xfer;
  --sysid_control_slave_in_a_read_cycle assignment, which is an e_assign
  sysid_control_slave_in_a_read_cycle <= ((internal_clock_crossing_0_m1_granted_sysid_control_slave AND clock_crossing_0_m1_read)) OR ((internal_clock_crossing_1_m1_granted_sysid_control_slave AND clock_crossing_1_m1_read));
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= sysid_control_slave_in_a_read_cycle;
  --sysid_control_slave_waits_for_write in a cycle, which is an e_mux
  sysid_control_slave_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(sysid_control_slave_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --sysid_control_slave_in_a_write_cycle assignment, which is an e_assign
  sysid_control_slave_in_a_write_cycle <= ((internal_clock_crossing_0_m1_granted_sysid_control_slave AND clock_crossing_0_m1_write)) OR ((internal_clock_crossing_1_m1_granted_sysid_control_slave AND clock_crossing_1_m1_write));
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= sysid_control_slave_in_a_write_cycle;
  wait_for_sysid_control_slave_counter <= std_logic'('0');
  --vhdl renameroo for output signals
  clock_crossing_0_m1_granted_sysid_control_slave <= internal_clock_crossing_0_m1_granted_sysid_control_slave;
  --vhdl renameroo for output signals
  clock_crossing_0_m1_qualified_request_sysid_control_slave <= internal_clock_crossing_0_m1_qualified_request_sysid_control_slave;
  --vhdl renameroo for output signals
  clock_crossing_0_m1_requests_sysid_control_slave <= internal_clock_crossing_0_m1_requests_sysid_control_slave;
  --vhdl renameroo for output signals
  clock_crossing_1_m1_granted_sysid_control_slave <= internal_clock_crossing_1_m1_granted_sysid_control_slave;
  --vhdl renameroo for output signals
  clock_crossing_1_m1_qualified_request_sysid_control_slave <= internal_clock_crossing_1_m1_qualified_request_sysid_control_slave;
  --vhdl renameroo for output signals
  clock_crossing_1_m1_requests_sysid_control_slave <= internal_clock_crossing_1_m1_requests_sysid_control_slave;
--synthesis translate_off
    --sysid/control_slave enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --grant signals are active simultaneously, which is an e_process
    process (clk)
    VARIABLE write_line49 : line;
    begin
      if clk'event and clk = '1' then
        if (std_logic_vector'("000000000000000000000000000000") & (((std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(internal_clock_crossing_0_m1_granted_sysid_control_slave))) + (std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(internal_clock_crossing_1_m1_granted_sysid_control_slave))))))>std_logic_vector'("00000000000000000000000000000001") then 
          write(write_line49, now);
          write(write_line49, string'(": "));
          write(write_line49, string'("> 1 of grant signals are active simultaneously"));
          write(output, write_line49.all);
          deallocate (write_line49);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --saved_grant signals are active simultaneously, which is an e_process
    process (clk)
    VARIABLE write_line50 : line;
    begin
      if clk'event and clk = '1' then
        if (std_logic_vector'("000000000000000000000000000000") & (((std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(clock_crossing_0_m1_saved_grant_sysid_control_slave))) + (std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(clock_crossing_1_m1_saved_grant_sysid_control_slave))))))>std_logic_vector'("00000000000000000000000000000001") then 
          write(write_line50, now);
          write(write_line50, string'(": "));
          write(write_line50, string'("> 1 of saved_grant signals are active simultaneously"));
          write(output, write_line50.all);
          deallocate (write_line50);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity system_timer_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal clock_crossing_0_m1_address_to_slave : IN STD_LOGIC_VECTOR (6 DOWNTO 0);
                 signal clock_crossing_0_m1_latency_counter : IN STD_LOGIC;
                 signal clock_crossing_0_m1_nativeaddress : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
                 signal clock_crossing_0_m1_read : IN STD_LOGIC;
                 signal clock_crossing_0_m1_write : IN STD_LOGIC;
                 signal clock_crossing_0_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;
                 signal system_timer_s1_irq : IN STD_LOGIC;
                 signal system_timer_s1_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

              -- outputs:
                 signal clock_crossing_0_m1_granted_system_timer_s1 : OUT STD_LOGIC;
                 signal clock_crossing_0_m1_qualified_request_system_timer_s1 : OUT STD_LOGIC;
                 signal clock_crossing_0_m1_read_data_valid_system_timer_s1 : OUT STD_LOGIC;
                 signal clock_crossing_0_m1_requests_system_timer_s1 : OUT STD_LOGIC;
                 signal d1_system_timer_s1_end_xfer : OUT STD_LOGIC;
                 signal system_timer_s1_address : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal system_timer_s1_chipselect : OUT STD_LOGIC;
                 signal system_timer_s1_irq_from_sa : OUT STD_LOGIC;
                 signal system_timer_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal system_timer_s1_reset_n : OUT STD_LOGIC;
                 signal system_timer_s1_write_n : OUT STD_LOGIC;
                 signal system_timer_s1_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
              );
end entity system_timer_s1_arbitrator;


architecture europa of system_timer_s1_arbitrator is
                signal clock_crossing_0_m1_arbiterlock :  STD_LOGIC;
                signal clock_crossing_0_m1_arbiterlock2 :  STD_LOGIC;
                signal clock_crossing_0_m1_continuerequest :  STD_LOGIC;
                signal clock_crossing_0_m1_saved_grant_system_timer_s1 :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_system_timer_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_clock_crossing_0_m1_granted_system_timer_s1 :  STD_LOGIC;
                signal internal_clock_crossing_0_m1_qualified_request_system_timer_s1 :  STD_LOGIC;
                signal internal_clock_crossing_0_m1_requests_system_timer_s1 :  STD_LOGIC;
                signal system_timer_s1_allgrants :  STD_LOGIC;
                signal system_timer_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal system_timer_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal system_timer_s1_any_continuerequest :  STD_LOGIC;
                signal system_timer_s1_arb_counter_enable :  STD_LOGIC;
                signal system_timer_s1_arb_share_counter :  STD_LOGIC;
                signal system_timer_s1_arb_share_counter_next_value :  STD_LOGIC;
                signal system_timer_s1_arb_share_set_values :  STD_LOGIC;
                signal system_timer_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal system_timer_s1_begins_xfer :  STD_LOGIC;
                signal system_timer_s1_end_xfer :  STD_LOGIC;
                signal system_timer_s1_firsttransfer :  STD_LOGIC;
                signal system_timer_s1_grant_vector :  STD_LOGIC;
                signal system_timer_s1_in_a_read_cycle :  STD_LOGIC;
                signal system_timer_s1_in_a_write_cycle :  STD_LOGIC;
                signal system_timer_s1_master_qreq_vector :  STD_LOGIC;
                signal system_timer_s1_non_bursting_master_requests :  STD_LOGIC;
                signal system_timer_s1_reg_firsttransfer :  STD_LOGIC;
                signal system_timer_s1_slavearbiterlockenable :  STD_LOGIC;
                signal system_timer_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal system_timer_s1_unreg_firsttransfer :  STD_LOGIC;
                signal system_timer_s1_waits_for_read :  STD_LOGIC;
                signal system_timer_s1_waits_for_write :  STD_LOGIC;
                signal wait_for_system_timer_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT system_timer_s1_end_xfer;
    end if;

  end process;

  system_timer_s1_begins_xfer <= NOT d1_reasons_to_wait AND (internal_clock_crossing_0_m1_qualified_request_system_timer_s1);
  --assign system_timer_s1_readdata_from_sa = system_timer_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  system_timer_s1_readdata_from_sa <= system_timer_s1_readdata;
  internal_clock_crossing_0_m1_requests_system_timer_s1 <= to_std_logic(((Std_Logic_Vector'(clock_crossing_0_m1_address_to_slave(6 DOWNTO 5) & std_logic_vector'("00000")) = std_logic_vector'("0000000")))) AND ((clock_crossing_0_m1_read OR clock_crossing_0_m1_write));
  --system_timer_s1_arb_share_counter set values, which is an e_mux
  system_timer_s1_arb_share_set_values <= std_logic'('1');
  --system_timer_s1_non_bursting_master_requests mux, which is an e_mux
  system_timer_s1_non_bursting_master_requests <= internal_clock_crossing_0_m1_requests_system_timer_s1;
  --system_timer_s1_any_bursting_master_saved_grant mux, which is an e_mux
  system_timer_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --system_timer_s1_arb_share_counter_next_value assignment, which is an e_assign
  system_timer_s1_arb_share_counter_next_value <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(system_timer_s1_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(system_timer_s1_arb_share_set_values))) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(system_timer_s1_arb_share_counter) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(system_timer_s1_arb_share_counter))) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))));
  --system_timer_s1_allgrants all slave grants, which is an e_mux
  system_timer_s1_allgrants <= system_timer_s1_grant_vector;
  --system_timer_s1_end_xfer assignment, which is an e_assign
  system_timer_s1_end_xfer <= NOT ((system_timer_s1_waits_for_read OR system_timer_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_system_timer_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_system_timer_s1 <= system_timer_s1_end_xfer AND (((NOT system_timer_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --system_timer_s1_arb_share_counter arbitration counter enable, which is an e_assign
  system_timer_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_system_timer_s1 AND system_timer_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_system_timer_s1 AND NOT system_timer_s1_non_bursting_master_requests));
  --system_timer_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      system_timer_s1_arb_share_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(system_timer_s1_arb_counter_enable) = '1' then 
        system_timer_s1_arb_share_counter <= system_timer_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --system_timer_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      system_timer_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((system_timer_s1_master_qreq_vector AND end_xfer_arb_share_counter_term_system_timer_s1)) OR ((end_xfer_arb_share_counter_term_system_timer_s1 AND NOT system_timer_s1_non_bursting_master_requests)))) = '1' then 
        system_timer_s1_slavearbiterlockenable <= system_timer_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --clock_crossing_0/m1 system_timer/s1 arbiterlock, which is an e_assign
  clock_crossing_0_m1_arbiterlock <= system_timer_s1_slavearbiterlockenable AND clock_crossing_0_m1_continuerequest;
  --system_timer_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  system_timer_s1_slavearbiterlockenable2 <= system_timer_s1_arb_share_counter_next_value;
  --clock_crossing_0/m1 system_timer/s1 arbiterlock2, which is an e_assign
  clock_crossing_0_m1_arbiterlock2 <= system_timer_s1_slavearbiterlockenable2 AND clock_crossing_0_m1_continuerequest;
  --system_timer_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  system_timer_s1_any_continuerequest <= std_logic'('1');
  --clock_crossing_0_m1_continuerequest continued request, which is an e_assign
  clock_crossing_0_m1_continuerequest <= std_logic'('1');
  internal_clock_crossing_0_m1_qualified_request_system_timer_s1 <= internal_clock_crossing_0_m1_requests_system_timer_s1 AND NOT ((clock_crossing_0_m1_read AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(clock_crossing_0_m1_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))))));
  --local readdatavalid clock_crossing_0_m1_read_data_valid_system_timer_s1, which is an e_mux
  clock_crossing_0_m1_read_data_valid_system_timer_s1 <= (internal_clock_crossing_0_m1_granted_system_timer_s1 AND clock_crossing_0_m1_read) AND NOT system_timer_s1_waits_for_read;
  --system_timer_s1_writedata mux, which is an e_mux
  system_timer_s1_writedata <= clock_crossing_0_m1_writedata (15 DOWNTO 0);
  --master is always granted when requested
  internal_clock_crossing_0_m1_granted_system_timer_s1 <= internal_clock_crossing_0_m1_qualified_request_system_timer_s1;
  --clock_crossing_0/m1 saved-grant system_timer/s1, which is an e_assign
  clock_crossing_0_m1_saved_grant_system_timer_s1 <= internal_clock_crossing_0_m1_requests_system_timer_s1;
  --allow new arb cycle for system_timer/s1, which is an e_assign
  system_timer_s1_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  system_timer_s1_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  system_timer_s1_master_qreq_vector <= std_logic'('1');
  --system_timer_s1_reset_n assignment, which is an e_assign
  system_timer_s1_reset_n <= reset_n;
  system_timer_s1_chipselect <= internal_clock_crossing_0_m1_granted_system_timer_s1;
  --system_timer_s1_firsttransfer first transaction, which is an e_assign
  system_timer_s1_firsttransfer <= A_WE_StdLogic((std_logic'(system_timer_s1_begins_xfer) = '1'), system_timer_s1_unreg_firsttransfer, system_timer_s1_reg_firsttransfer);
  --system_timer_s1_unreg_firsttransfer first transaction, which is an e_assign
  system_timer_s1_unreg_firsttransfer <= NOT ((system_timer_s1_slavearbiterlockenable AND system_timer_s1_any_continuerequest));
  --system_timer_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      system_timer_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(system_timer_s1_begins_xfer) = '1' then 
        system_timer_s1_reg_firsttransfer <= system_timer_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --system_timer_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  system_timer_s1_beginbursttransfer_internal <= system_timer_s1_begins_xfer;
  --~system_timer_s1_write_n assignment, which is an e_mux
  system_timer_s1_write_n <= NOT ((internal_clock_crossing_0_m1_granted_system_timer_s1 AND clock_crossing_0_m1_write));
  --system_timer_s1_address mux, which is an e_mux
  system_timer_s1_address <= clock_crossing_0_m1_nativeaddress (2 DOWNTO 0);
  --d1_system_timer_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_system_timer_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_system_timer_s1_end_xfer <= system_timer_s1_end_xfer;
    end if;

  end process;

  --system_timer_s1_waits_for_read in a cycle, which is an e_mux
  system_timer_s1_waits_for_read <= system_timer_s1_in_a_read_cycle AND system_timer_s1_begins_xfer;
  --system_timer_s1_in_a_read_cycle assignment, which is an e_assign
  system_timer_s1_in_a_read_cycle <= internal_clock_crossing_0_m1_granted_system_timer_s1 AND clock_crossing_0_m1_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= system_timer_s1_in_a_read_cycle;
  --system_timer_s1_waits_for_write in a cycle, which is an e_mux
  system_timer_s1_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(system_timer_s1_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --system_timer_s1_in_a_write_cycle assignment, which is an e_assign
  system_timer_s1_in_a_write_cycle <= internal_clock_crossing_0_m1_granted_system_timer_s1 AND clock_crossing_0_m1_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= system_timer_s1_in_a_write_cycle;
  wait_for_system_timer_s1_counter <= std_logic'('0');
  --assign system_timer_s1_irq_from_sa = system_timer_s1_irq so that symbol knows where to group signals which may go to master only, which is an e_assign
  system_timer_s1_irq_from_sa <= system_timer_s1_irq;
  --vhdl renameroo for output signals
  clock_crossing_0_m1_granted_system_timer_s1 <= internal_clock_crossing_0_m1_granted_system_timer_s1;
  --vhdl renameroo for output signals
  clock_crossing_0_m1_qualified_request_system_timer_s1 <= internal_clock_crossing_0_m1_qualified_request_system_timer_s1;
  --vhdl renameroo for output signals
  clock_crossing_0_m1_requests_system_timer_s1 <= internal_clock_crossing_0_m1_requests_system_timer_s1;
--synthesis translate_off
    --system_timer/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity system_timer_ap_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal clock_crossing_1_m1_address_to_slave : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal clock_crossing_1_m1_latency_counter : IN STD_LOGIC;
                 signal clock_crossing_1_m1_nativeaddress : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
                 signal clock_crossing_1_m1_read : IN STD_LOGIC;
                 signal clock_crossing_1_m1_write : IN STD_LOGIC;
                 signal clock_crossing_1_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;
                 signal system_timer_ap_s1_irq : IN STD_LOGIC;
                 signal system_timer_ap_s1_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

              -- outputs:
                 signal clock_crossing_1_m1_granted_system_timer_ap_s1 : OUT STD_LOGIC;
                 signal clock_crossing_1_m1_qualified_request_system_timer_ap_s1 : OUT STD_LOGIC;
                 signal clock_crossing_1_m1_read_data_valid_system_timer_ap_s1 : OUT STD_LOGIC;
                 signal clock_crossing_1_m1_requests_system_timer_ap_s1 : OUT STD_LOGIC;
                 signal d1_system_timer_ap_s1_end_xfer : OUT STD_LOGIC;
                 signal system_timer_ap_s1_address : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal system_timer_ap_s1_chipselect : OUT STD_LOGIC;
                 signal system_timer_ap_s1_irq_from_sa : OUT STD_LOGIC;
                 signal system_timer_ap_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal system_timer_ap_s1_reset_n : OUT STD_LOGIC;
                 signal system_timer_ap_s1_write_n : OUT STD_LOGIC;
                 signal system_timer_ap_s1_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
              );
end entity system_timer_ap_s1_arbitrator;


architecture europa of system_timer_ap_s1_arbitrator is
                signal clock_crossing_1_m1_arbiterlock :  STD_LOGIC;
                signal clock_crossing_1_m1_arbiterlock2 :  STD_LOGIC;
                signal clock_crossing_1_m1_continuerequest :  STD_LOGIC;
                signal clock_crossing_1_m1_saved_grant_system_timer_ap_s1 :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_system_timer_ap_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_clock_crossing_1_m1_granted_system_timer_ap_s1 :  STD_LOGIC;
                signal internal_clock_crossing_1_m1_qualified_request_system_timer_ap_s1 :  STD_LOGIC;
                signal internal_clock_crossing_1_m1_requests_system_timer_ap_s1 :  STD_LOGIC;
                signal system_timer_ap_s1_allgrants :  STD_LOGIC;
                signal system_timer_ap_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal system_timer_ap_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal system_timer_ap_s1_any_continuerequest :  STD_LOGIC;
                signal system_timer_ap_s1_arb_counter_enable :  STD_LOGIC;
                signal system_timer_ap_s1_arb_share_counter :  STD_LOGIC;
                signal system_timer_ap_s1_arb_share_counter_next_value :  STD_LOGIC;
                signal system_timer_ap_s1_arb_share_set_values :  STD_LOGIC;
                signal system_timer_ap_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal system_timer_ap_s1_begins_xfer :  STD_LOGIC;
                signal system_timer_ap_s1_end_xfer :  STD_LOGIC;
                signal system_timer_ap_s1_firsttransfer :  STD_LOGIC;
                signal system_timer_ap_s1_grant_vector :  STD_LOGIC;
                signal system_timer_ap_s1_in_a_read_cycle :  STD_LOGIC;
                signal system_timer_ap_s1_in_a_write_cycle :  STD_LOGIC;
                signal system_timer_ap_s1_master_qreq_vector :  STD_LOGIC;
                signal system_timer_ap_s1_non_bursting_master_requests :  STD_LOGIC;
                signal system_timer_ap_s1_reg_firsttransfer :  STD_LOGIC;
                signal system_timer_ap_s1_slavearbiterlockenable :  STD_LOGIC;
                signal system_timer_ap_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal system_timer_ap_s1_unreg_firsttransfer :  STD_LOGIC;
                signal system_timer_ap_s1_waits_for_read :  STD_LOGIC;
                signal system_timer_ap_s1_waits_for_write :  STD_LOGIC;
                signal wait_for_system_timer_ap_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT system_timer_ap_s1_end_xfer;
    end if;

  end process;

  system_timer_ap_s1_begins_xfer <= NOT d1_reasons_to_wait AND (internal_clock_crossing_1_m1_qualified_request_system_timer_ap_s1);
  --assign system_timer_ap_s1_readdata_from_sa = system_timer_ap_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  system_timer_ap_s1_readdata_from_sa <= system_timer_ap_s1_readdata;
  internal_clock_crossing_1_m1_requests_system_timer_ap_s1 <= to_std_logic(((Std_Logic_Vector'(clock_crossing_1_m1_address_to_slave(7 DOWNTO 5) & std_logic_vector'("00000")) = std_logic_vector'("10000000")))) AND ((clock_crossing_1_m1_read OR clock_crossing_1_m1_write));
  --system_timer_ap_s1_arb_share_counter set values, which is an e_mux
  system_timer_ap_s1_arb_share_set_values <= std_logic'('1');
  --system_timer_ap_s1_non_bursting_master_requests mux, which is an e_mux
  system_timer_ap_s1_non_bursting_master_requests <= internal_clock_crossing_1_m1_requests_system_timer_ap_s1;
  --system_timer_ap_s1_any_bursting_master_saved_grant mux, which is an e_mux
  system_timer_ap_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --system_timer_ap_s1_arb_share_counter_next_value assignment, which is an e_assign
  system_timer_ap_s1_arb_share_counter_next_value <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(system_timer_ap_s1_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(system_timer_ap_s1_arb_share_set_values))) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(system_timer_ap_s1_arb_share_counter) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(system_timer_ap_s1_arb_share_counter))) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))));
  --system_timer_ap_s1_allgrants all slave grants, which is an e_mux
  system_timer_ap_s1_allgrants <= system_timer_ap_s1_grant_vector;
  --system_timer_ap_s1_end_xfer assignment, which is an e_assign
  system_timer_ap_s1_end_xfer <= NOT ((system_timer_ap_s1_waits_for_read OR system_timer_ap_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_system_timer_ap_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_system_timer_ap_s1 <= system_timer_ap_s1_end_xfer AND (((NOT system_timer_ap_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --system_timer_ap_s1_arb_share_counter arbitration counter enable, which is an e_assign
  system_timer_ap_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_system_timer_ap_s1 AND system_timer_ap_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_system_timer_ap_s1 AND NOT system_timer_ap_s1_non_bursting_master_requests));
  --system_timer_ap_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      system_timer_ap_s1_arb_share_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(system_timer_ap_s1_arb_counter_enable) = '1' then 
        system_timer_ap_s1_arb_share_counter <= system_timer_ap_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --system_timer_ap_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      system_timer_ap_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((system_timer_ap_s1_master_qreq_vector AND end_xfer_arb_share_counter_term_system_timer_ap_s1)) OR ((end_xfer_arb_share_counter_term_system_timer_ap_s1 AND NOT system_timer_ap_s1_non_bursting_master_requests)))) = '1' then 
        system_timer_ap_s1_slavearbiterlockenable <= system_timer_ap_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --clock_crossing_1/m1 system_timer_ap/s1 arbiterlock, which is an e_assign
  clock_crossing_1_m1_arbiterlock <= system_timer_ap_s1_slavearbiterlockenable AND clock_crossing_1_m1_continuerequest;
  --system_timer_ap_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  system_timer_ap_s1_slavearbiterlockenable2 <= system_timer_ap_s1_arb_share_counter_next_value;
  --clock_crossing_1/m1 system_timer_ap/s1 arbiterlock2, which is an e_assign
  clock_crossing_1_m1_arbiterlock2 <= system_timer_ap_s1_slavearbiterlockenable2 AND clock_crossing_1_m1_continuerequest;
  --system_timer_ap_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  system_timer_ap_s1_any_continuerequest <= std_logic'('1');
  --clock_crossing_1_m1_continuerequest continued request, which is an e_assign
  clock_crossing_1_m1_continuerequest <= std_logic'('1');
  internal_clock_crossing_1_m1_qualified_request_system_timer_ap_s1 <= internal_clock_crossing_1_m1_requests_system_timer_ap_s1 AND NOT ((clock_crossing_1_m1_read AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(clock_crossing_1_m1_latency_counter))) /= std_logic_vector'("00000000000000000000000000000000"))))));
  --local readdatavalid clock_crossing_1_m1_read_data_valid_system_timer_ap_s1, which is an e_mux
  clock_crossing_1_m1_read_data_valid_system_timer_ap_s1 <= (internal_clock_crossing_1_m1_granted_system_timer_ap_s1 AND clock_crossing_1_m1_read) AND NOT system_timer_ap_s1_waits_for_read;
  --system_timer_ap_s1_writedata mux, which is an e_mux
  system_timer_ap_s1_writedata <= clock_crossing_1_m1_writedata (15 DOWNTO 0);
  --master is always granted when requested
  internal_clock_crossing_1_m1_granted_system_timer_ap_s1 <= internal_clock_crossing_1_m1_qualified_request_system_timer_ap_s1;
  --clock_crossing_1/m1 saved-grant system_timer_ap/s1, which is an e_assign
  clock_crossing_1_m1_saved_grant_system_timer_ap_s1 <= internal_clock_crossing_1_m1_requests_system_timer_ap_s1;
  --allow new arb cycle for system_timer_ap/s1, which is an e_assign
  system_timer_ap_s1_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  system_timer_ap_s1_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  system_timer_ap_s1_master_qreq_vector <= std_logic'('1');
  --system_timer_ap_s1_reset_n assignment, which is an e_assign
  system_timer_ap_s1_reset_n <= reset_n;
  system_timer_ap_s1_chipselect <= internal_clock_crossing_1_m1_granted_system_timer_ap_s1;
  --system_timer_ap_s1_firsttransfer first transaction, which is an e_assign
  system_timer_ap_s1_firsttransfer <= A_WE_StdLogic((std_logic'(system_timer_ap_s1_begins_xfer) = '1'), system_timer_ap_s1_unreg_firsttransfer, system_timer_ap_s1_reg_firsttransfer);
  --system_timer_ap_s1_unreg_firsttransfer first transaction, which is an e_assign
  system_timer_ap_s1_unreg_firsttransfer <= NOT ((system_timer_ap_s1_slavearbiterlockenable AND system_timer_ap_s1_any_continuerequest));
  --system_timer_ap_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      system_timer_ap_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(system_timer_ap_s1_begins_xfer) = '1' then 
        system_timer_ap_s1_reg_firsttransfer <= system_timer_ap_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --system_timer_ap_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  system_timer_ap_s1_beginbursttransfer_internal <= system_timer_ap_s1_begins_xfer;
  --~system_timer_ap_s1_write_n assignment, which is an e_mux
  system_timer_ap_s1_write_n <= NOT ((internal_clock_crossing_1_m1_granted_system_timer_ap_s1 AND clock_crossing_1_m1_write));
  --system_timer_ap_s1_address mux, which is an e_mux
  system_timer_ap_s1_address <= clock_crossing_1_m1_nativeaddress (2 DOWNTO 0);
  --d1_system_timer_ap_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_system_timer_ap_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_system_timer_ap_s1_end_xfer <= system_timer_ap_s1_end_xfer;
    end if;

  end process;

  --system_timer_ap_s1_waits_for_read in a cycle, which is an e_mux
  system_timer_ap_s1_waits_for_read <= system_timer_ap_s1_in_a_read_cycle AND system_timer_ap_s1_begins_xfer;
  --system_timer_ap_s1_in_a_read_cycle assignment, which is an e_assign
  system_timer_ap_s1_in_a_read_cycle <= internal_clock_crossing_1_m1_granted_system_timer_ap_s1 AND clock_crossing_1_m1_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= system_timer_ap_s1_in_a_read_cycle;
  --system_timer_ap_s1_waits_for_write in a cycle, which is an e_mux
  system_timer_ap_s1_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(system_timer_ap_s1_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --system_timer_ap_s1_in_a_write_cycle assignment, which is an e_assign
  system_timer_ap_s1_in_a_write_cycle <= internal_clock_crossing_1_m1_granted_system_timer_ap_s1 AND clock_crossing_1_m1_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= system_timer_ap_s1_in_a_write_cycle;
  wait_for_system_timer_ap_s1_counter <= std_logic'('0');
  --assign system_timer_ap_s1_irq_from_sa = system_timer_ap_s1_irq so that symbol knows where to group signals which may go to master only, which is an e_assign
  system_timer_ap_s1_irq_from_sa <= system_timer_ap_s1_irq;
  --vhdl renameroo for output signals
  clock_crossing_1_m1_granted_system_timer_ap_s1 <= internal_clock_crossing_1_m1_granted_system_timer_ap_s1;
  --vhdl renameroo for output signals
  clock_crossing_1_m1_qualified_request_system_timer_ap_s1 <= internal_clock_crossing_1_m1_qualified_request_system_timer_ap_s1;
  --vhdl renameroo for output signals
  clock_crossing_1_m1_requests_system_timer_ap_s1 <= internal_clock_crossing_1_m1_requests_system_timer_ap_s1;
--synthesis translate_off
    --system_timer_ap/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity tri_state_bridge_0_avalon_slave_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal pcp_cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (25 DOWNTO 0);
                 signal pcp_cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal pcp_cpu_data_master_dbs_address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal pcp_cpu_data_master_dbs_write_16 : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal pcp_cpu_data_master_no_byte_enables_and_last_term : IN STD_LOGIC;
                 signal pcp_cpu_data_master_read : IN STD_LOGIC;
                 signal pcp_cpu_data_master_write : IN STD_LOGIC;
                 signal pcp_cpu_instruction_master_address_to_slave : IN STD_LOGIC_VECTOR (25 DOWNTO 0);
                 signal pcp_cpu_instruction_master_dbs_address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal pcp_cpu_instruction_master_latency_counter : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal pcp_cpu_instruction_master_read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal DBC3C40_SRAM_0_avalon_tristate_slave_wait_counter_eq_0 : OUT STD_LOGIC;
                 signal ben_to_the_DBC3C40_SRAM_0 : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal cfi_flash_0_s1_wait_counter_eq_0 : OUT STD_LOGIC;
                 signal cfi_flash_0_s1_wait_counter_eq_1 : OUT STD_LOGIC;
                 signal d1_tri_state_bridge_0_avalon_slave_end_xfer : OUT STD_LOGIC;
                 signal incoming_tri_state_bridge_0_data : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal incoming_tri_state_bridge_0_data_with_Xs_converted_to_0 : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal ncs_to_the_DBC3C40_SRAM_0 : OUT STD_LOGIC;
                 signal pcp_cpu_data_master_byteenable_DBC3C40_SRAM_0_avalon_tristate_slave : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal pcp_cpu_data_master_byteenable_cfi_flash_0_s1 : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal pcp_cpu_data_master_granted_DBC3C40_SRAM_0_avalon_tristate_slave : OUT STD_LOGIC;
                 signal pcp_cpu_data_master_granted_cfi_flash_0_s1 : OUT STD_LOGIC;
                 signal pcp_cpu_data_master_qualified_request_DBC3C40_SRAM_0_avalon_tristate_slave : OUT STD_LOGIC;
                 signal pcp_cpu_data_master_qualified_request_cfi_flash_0_s1 : OUT STD_LOGIC;
                 signal pcp_cpu_data_master_read_data_valid_DBC3C40_SRAM_0_avalon_tristate_slave : OUT STD_LOGIC;
                 signal pcp_cpu_data_master_read_data_valid_cfi_flash_0_s1 : OUT STD_LOGIC;
                 signal pcp_cpu_data_master_requests_DBC3C40_SRAM_0_avalon_tristate_slave : OUT STD_LOGIC;
                 signal pcp_cpu_data_master_requests_cfi_flash_0_s1 : OUT STD_LOGIC;
                 signal pcp_cpu_instruction_master_granted_DBC3C40_SRAM_0_avalon_tristate_slave : OUT STD_LOGIC;
                 signal pcp_cpu_instruction_master_granted_cfi_flash_0_s1 : OUT STD_LOGIC;
                 signal pcp_cpu_instruction_master_qualified_request_DBC3C40_SRAM_0_avalon_tristate_slave : OUT STD_LOGIC;
                 signal pcp_cpu_instruction_master_qualified_request_cfi_flash_0_s1 : OUT STD_LOGIC;
                 signal pcp_cpu_instruction_master_read_data_valid_DBC3C40_SRAM_0_avalon_tristate_slave : OUT STD_LOGIC;
                 signal pcp_cpu_instruction_master_read_data_valid_cfi_flash_0_s1 : OUT STD_LOGIC;
                 signal pcp_cpu_instruction_master_requests_DBC3C40_SRAM_0_avalon_tristate_slave : OUT STD_LOGIC;
                 signal pcp_cpu_instruction_master_requests_cfi_flash_0_s1 : OUT STD_LOGIC;
                 signal registered_pcp_cpu_data_master_read_data_valid_DBC3C40_SRAM_0_avalon_tristate_slave : OUT STD_LOGIC;
                 signal registered_pcp_cpu_data_master_read_data_valid_cfi_flash_0_s1 : OUT STD_LOGIC;
                 signal select_n_to_the_cfi_flash_0 : OUT STD_LOGIC;
                 signal tri_state_bridge_0_address : OUT STD_LOGIC_VECTOR (22 DOWNTO 0);
                 signal tri_state_bridge_0_data : INOUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal tri_state_bridge_0_readn : OUT STD_LOGIC;
                 signal tri_state_bridge_0_writen : OUT STD_LOGIC
              );
end entity tri_state_bridge_0_avalon_slave_arbitrator;


architecture europa of tri_state_bridge_0_avalon_slave_arbitrator is
                signal DBC3C40_SRAM_0_avalon_tristate_slave_counter_load_value :  STD_LOGIC;
                signal DBC3C40_SRAM_0_avalon_tristate_slave_in_a_read_cycle :  STD_LOGIC;
                signal DBC3C40_SRAM_0_avalon_tristate_slave_in_a_write_cycle :  STD_LOGIC;
                signal DBC3C40_SRAM_0_avalon_tristate_slave_wait_counter :  STD_LOGIC;
                signal DBC3C40_SRAM_0_avalon_tristate_slave_waits_for_read :  STD_LOGIC;
                signal DBC3C40_SRAM_0_avalon_tristate_slave_waits_for_write :  STD_LOGIC;
                signal DBC3C40_SRAM_0_avalon_tristate_slave_with_write_latency :  STD_LOGIC;
                signal cfi_flash_0_s1_counter_load_value :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal cfi_flash_0_s1_in_a_read_cycle :  STD_LOGIC;
                signal cfi_flash_0_s1_in_a_write_cycle :  STD_LOGIC;
                signal cfi_flash_0_s1_wait_counter :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal cfi_flash_0_s1_waits_for_read :  STD_LOGIC;
                signal cfi_flash_0_s1_waits_for_write :  STD_LOGIC;
                signal cfi_flash_0_s1_with_write_latency :  STD_LOGIC;
                signal d1_in_a_write_cycle :  STD_LOGIC;
                signal d1_outgoing_tri_state_bridge_0_data :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_tri_state_bridge_0_avalon_slave :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal incoming_tri_state_bridge_0_data_bit_0_is_x :  STD_LOGIC;
                signal incoming_tri_state_bridge_0_data_bit_10_is_x :  STD_LOGIC;
                signal incoming_tri_state_bridge_0_data_bit_11_is_x :  STD_LOGIC;
                signal incoming_tri_state_bridge_0_data_bit_12_is_x :  STD_LOGIC;
                signal incoming_tri_state_bridge_0_data_bit_13_is_x :  STD_LOGIC;
                signal incoming_tri_state_bridge_0_data_bit_14_is_x :  STD_LOGIC;
                signal incoming_tri_state_bridge_0_data_bit_15_is_x :  STD_LOGIC;
                signal incoming_tri_state_bridge_0_data_bit_1_is_x :  STD_LOGIC;
                signal incoming_tri_state_bridge_0_data_bit_2_is_x :  STD_LOGIC;
                signal incoming_tri_state_bridge_0_data_bit_3_is_x :  STD_LOGIC;
                signal incoming_tri_state_bridge_0_data_bit_4_is_x :  STD_LOGIC;
                signal incoming_tri_state_bridge_0_data_bit_5_is_x :  STD_LOGIC;
                signal incoming_tri_state_bridge_0_data_bit_6_is_x :  STD_LOGIC;
                signal incoming_tri_state_bridge_0_data_bit_7_is_x :  STD_LOGIC;
                signal incoming_tri_state_bridge_0_data_bit_8_is_x :  STD_LOGIC;
                signal incoming_tri_state_bridge_0_data_bit_9_is_x :  STD_LOGIC;
                signal internal_DBC3C40_SRAM_0_avalon_tristate_slave_wait_counter_eq_0 :  STD_LOGIC;
                signal internal_cfi_flash_0_s1_wait_counter_eq_0 :  STD_LOGIC;
                signal internal_incoming_tri_state_bridge_0_data :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal internal_pcp_cpu_data_master_byteenable_DBC3C40_SRAM_0_avalon_tristate_slave :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal internal_pcp_cpu_data_master_byteenable_cfi_flash_0_s1 :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal internal_pcp_cpu_data_master_granted_DBC3C40_SRAM_0_avalon_tristate_slave :  STD_LOGIC;
                signal internal_pcp_cpu_data_master_granted_cfi_flash_0_s1 :  STD_LOGIC;
                signal internal_pcp_cpu_data_master_qualified_request_DBC3C40_SRAM_0_avalon_tristate_slave :  STD_LOGIC;
                signal internal_pcp_cpu_data_master_qualified_request_cfi_flash_0_s1 :  STD_LOGIC;
                signal internal_pcp_cpu_data_master_requests_DBC3C40_SRAM_0_avalon_tristate_slave :  STD_LOGIC;
                signal internal_pcp_cpu_data_master_requests_cfi_flash_0_s1 :  STD_LOGIC;
                signal internal_pcp_cpu_instruction_master_granted_DBC3C40_SRAM_0_avalon_tristate_slave :  STD_LOGIC;
                signal internal_pcp_cpu_instruction_master_granted_cfi_flash_0_s1 :  STD_LOGIC;
                signal internal_pcp_cpu_instruction_master_qualified_request_DBC3C40_SRAM_0_avalon_tristate_slave :  STD_LOGIC;
                signal internal_pcp_cpu_instruction_master_qualified_request_cfi_flash_0_s1 :  STD_LOGIC;
                signal internal_pcp_cpu_instruction_master_requests_DBC3C40_SRAM_0_avalon_tristate_slave :  STD_LOGIC;
                signal internal_pcp_cpu_instruction_master_requests_cfi_flash_0_s1 :  STD_LOGIC;
                signal last_cycle_pcp_cpu_data_master_granted_slave_DBC3C40_SRAM_0_avalon_tristate_slave :  STD_LOGIC;
                signal last_cycle_pcp_cpu_data_master_granted_slave_cfi_flash_0_s1 :  STD_LOGIC;
                signal last_cycle_pcp_cpu_instruction_master_granted_slave_DBC3C40_SRAM_0_avalon_tristate_slave :  STD_LOGIC;
                signal last_cycle_pcp_cpu_instruction_master_granted_slave_cfi_flash_0_s1 :  STD_LOGIC;
                signal outgoing_tri_state_bridge_0_data :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal p1_ben_to_the_DBC3C40_SRAM_0 :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal p1_ncs_to_the_DBC3C40_SRAM_0 :  STD_LOGIC;
                signal p1_pcp_cpu_data_master_read_data_valid_DBC3C40_SRAM_0_avalon_tristate_slave_shift_register :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal p1_pcp_cpu_data_master_read_data_valid_cfi_flash_0_s1_shift_register :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal p1_pcp_cpu_instruction_master_read_data_valid_DBC3C40_SRAM_0_avalon_tristate_slave_shift_register :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal p1_pcp_cpu_instruction_master_read_data_valid_cfi_flash_0_s1_shift_register :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal p1_select_n_to_the_cfi_flash_0 :  STD_LOGIC;
                signal p1_tri_state_bridge_0_address :  STD_LOGIC_VECTOR (22 DOWNTO 0);
                signal p1_tri_state_bridge_0_readn :  STD_LOGIC;
                signal p1_tri_state_bridge_0_writen :  STD_LOGIC;
                signal pcp_cpu_data_master_arbiterlock :  STD_LOGIC;
                signal pcp_cpu_data_master_arbiterlock2 :  STD_LOGIC;
                signal pcp_cpu_data_master_byteenable_DBC3C40_SRAM_0_avalon_tristate_slave_segment_0 :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal pcp_cpu_data_master_byteenable_DBC3C40_SRAM_0_avalon_tristate_slave_segment_1 :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal pcp_cpu_data_master_byteenable_cfi_flash_0_s1_segment_0 :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal pcp_cpu_data_master_byteenable_cfi_flash_0_s1_segment_1 :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal pcp_cpu_data_master_continuerequest :  STD_LOGIC;
                signal pcp_cpu_data_master_read_data_valid_DBC3C40_SRAM_0_avalon_tristate_slave_shift_register :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal pcp_cpu_data_master_read_data_valid_DBC3C40_SRAM_0_avalon_tristate_slave_shift_register_in :  STD_LOGIC;
                signal pcp_cpu_data_master_read_data_valid_cfi_flash_0_s1_shift_register :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal pcp_cpu_data_master_read_data_valid_cfi_flash_0_s1_shift_register_in :  STD_LOGIC;
                signal pcp_cpu_data_master_saved_grant_DBC3C40_SRAM_0_avalon_tristate_slave :  STD_LOGIC;
                signal pcp_cpu_data_master_saved_grant_cfi_flash_0_s1 :  STD_LOGIC;
                signal pcp_cpu_instruction_master_arbiterlock :  STD_LOGIC;
                signal pcp_cpu_instruction_master_arbiterlock2 :  STD_LOGIC;
                signal pcp_cpu_instruction_master_continuerequest :  STD_LOGIC;
                signal pcp_cpu_instruction_master_read_data_valid_DBC3C40_SRAM_0_avalon_tristate_slave_shift_register :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal pcp_cpu_instruction_master_read_data_valid_DBC3C40_SRAM_0_avalon_tristate_slave_shift_register_in :  STD_LOGIC;
                signal pcp_cpu_instruction_master_read_data_valid_cfi_flash_0_s1_shift_register :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal pcp_cpu_instruction_master_read_data_valid_cfi_flash_0_s1_shift_register_in :  STD_LOGIC;
                signal pcp_cpu_instruction_master_saved_grant_DBC3C40_SRAM_0_avalon_tristate_slave :  STD_LOGIC;
                signal pcp_cpu_instruction_master_saved_grant_cfi_flash_0_s1 :  STD_LOGIC;
                signal time_to_write :  STD_LOGIC;
                signal tri_state_bridge_0_avalon_slave_allgrants :  STD_LOGIC;
                signal tri_state_bridge_0_avalon_slave_allow_new_arb_cycle :  STD_LOGIC;
                signal tri_state_bridge_0_avalon_slave_any_bursting_master_saved_grant :  STD_LOGIC;
                signal tri_state_bridge_0_avalon_slave_any_continuerequest :  STD_LOGIC;
                signal tri_state_bridge_0_avalon_slave_arb_addend :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal tri_state_bridge_0_avalon_slave_arb_counter_enable :  STD_LOGIC;
                signal tri_state_bridge_0_avalon_slave_arb_share_counter :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal tri_state_bridge_0_avalon_slave_arb_share_counter_next_value :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal tri_state_bridge_0_avalon_slave_arb_share_set_values :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal tri_state_bridge_0_avalon_slave_arb_winner :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal tri_state_bridge_0_avalon_slave_arbitration_holdoff_internal :  STD_LOGIC;
                signal tri_state_bridge_0_avalon_slave_beginbursttransfer_internal :  STD_LOGIC;
                signal tri_state_bridge_0_avalon_slave_begins_xfer :  STD_LOGIC;
                signal tri_state_bridge_0_avalon_slave_chosen_master_double_vector :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal tri_state_bridge_0_avalon_slave_chosen_master_rot_left :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal tri_state_bridge_0_avalon_slave_end_xfer :  STD_LOGIC;
                signal tri_state_bridge_0_avalon_slave_firsttransfer :  STD_LOGIC;
                signal tri_state_bridge_0_avalon_slave_grant_vector :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal tri_state_bridge_0_avalon_slave_master_qreq_vector :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal tri_state_bridge_0_avalon_slave_non_bursting_master_requests :  STD_LOGIC;
                signal tri_state_bridge_0_avalon_slave_read_pending :  STD_LOGIC;
                signal tri_state_bridge_0_avalon_slave_reg_firsttransfer :  STD_LOGIC;
                signal tri_state_bridge_0_avalon_slave_saved_chosen_master_vector :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal tri_state_bridge_0_avalon_slave_slavearbiterlockenable :  STD_LOGIC;
                signal tri_state_bridge_0_avalon_slave_slavearbiterlockenable2 :  STD_LOGIC;
                signal tri_state_bridge_0_avalon_slave_unreg_firsttransfer :  STD_LOGIC;
                signal tri_state_bridge_0_avalon_slave_write_pending :  STD_LOGIC;
                signal wait_for_DBC3C40_SRAM_0_avalon_tristate_slave_counter :  STD_LOGIC;
                signal wait_for_cfi_flash_0_s1_counter :  STD_LOGIC;
attribute ALTERA_ATTRIBUTE : string;
attribute ALTERA_ATTRIBUTE of ben_to_the_DBC3C40_SRAM_0 : signal is "FAST_OUTPUT_REGISTER=ON";
attribute ALTERA_ATTRIBUTE of d1_in_a_write_cycle : signal is "FAST_OUTPUT_ENABLE_REGISTER=ON";
attribute ALTERA_ATTRIBUTE of d1_outgoing_tri_state_bridge_0_data : signal is "FAST_OUTPUT_REGISTER=ON";
attribute ALTERA_ATTRIBUTE of internal_incoming_tri_state_bridge_0_data : signal is "FAST_INPUT_REGISTER=ON";
attribute ALTERA_ATTRIBUTE of ncs_to_the_DBC3C40_SRAM_0 : signal is "FAST_OUTPUT_REGISTER=ON";
attribute ALTERA_ATTRIBUTE of select_n_to_the_cfi_flash_0 : signal is "FAST_OUTPUT_REGISTER=ON";
attribute ALTERA_ATTRIBUTE of tri_state_bridge_0_address : signal is "FAST_OUTPUT_REGISTER=ON";
attribute ALTERA_ATTRIBUTE of tri_state_bridge_0_readn : signal is "FAST_OUTPUT_REGISTER=ON";
attribute ALTERA_ATTRIBUTE of tri_state_bridge_0_writen : signal is "FAST_OUTPUT_REGISTER=ON";

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT tri_state_bridge_0_avalon_slave_end_xfer;
    end if;

  end process;

  tri_state_bridge_0_avalon_slave_begins_xfer <= NOT d1_reasons_to_wait AND ((((internal_pcp_cpu_data_master_qualified_request_DBC3C40_SRAM_0_avalon_tristate_slave OR internal_pcp_cpu_instruction_master_qualified_request_DBC3C40_SRAM_0_avalon_tristate_slave) OR internal_pcp_cpu_data_master_qualified_request_cfi_flash_0_s1) OR internal_pcp_cpu_instruction_master_qualified_request_cfi_flash_0_s1));
  internal_pcp_cpu_data_master_requests_DBC3C40_SRAM_0_avalon_tristate_slave <= to_std_logic(((Std_Logic_Vector'(pcp_cpu_data_master_address_to_slave(25 DOWNTO 20) & std_logic_vector'("00000000000000000000")) = std_logic_vector'("00001000000000000000000000")))) AND ((pcp_cpu_data_master_read OR pcp_cpu_data_master_write));
  --~ncs_to_the_DBC3C40_SRAM_0 of type chipselect to ~p1_ncs_to_the_DBC3C40_SRAM_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      ncs_to_the_DBC3C40_SRAM_0 <= Vector_To_Std_Logic(NOT std_logic_vector'("00000000000000000000000000000000"));
    elsif clk'event and clk = '1' then
      ncs_to_the_DBC3C40_SRAM_0 <= p1_ncs_to_the_DBC3C40_SRAM_0;
    end if;

  end process;

  --~select_n_to_the_cfi_flash_0 of type chipselect to ~p1_select_n_to_the_cfi_flash_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      select_n_to_the_cfi_flash_0 <= Vector_To_Std_Logic(NOT std_logic_vector'("00000000000000000000000000000000"));
    elsif clk'event and clk = '1' then
      select_n_to_the_cfi_flash_0 <= p1_select_n_to_the_cfi_flash_0;
    end if;

  end process;

  tri_state_bridge_0_avalon_slave_write_pending <= std_logic'('0');
  --tri_state_bridge_0/avalon_slave read pending calc, which is an e_assign
  tri_state_bridge_0_avalon_slave_read_pending <= std_logic'('0');
  --registered rdv signal_name registered_pcp_cpu_data_master_read_data_valid_DBC3C40_SRAM_0_avalon_tristate_slave assignment, which is an e_assign
  registered_pcp_cpu_data_master_read_data_valid_DBC3C40_SRAM_0_avalon_tristate_slave <= pcp_cpu_data_master_read_data_valid_DBC3C40_SRAM_0_avalon_tristate_slave_shift_register(0);
  --tri_state_bridge_0_avalon_slave_arb_share_counter set values, which is an e_mux
  tri_state_bridge_0_avalon_slave_arb_share_set_values <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_pcp_cpu_data_master_granted_DBC3C40_SRAM_0_avalon_tristate_slave)) = '1'), std_logic_vector'("00000000000000000000000000000010"), A_WE_StdLogicVector((std_logic'((internal_pcp_cpu_instruction_master_granted_DBC3C40_SRAM_0_avalon_tristate_slave)) = '1'), std_logic_vector'("00000000000000000000000000000010"), A_WE_StdLogicVector((std_logic'((internal_pcp_cpu_data_master_granted_cfi_flash_0_s1)) = '1'), std_logic_vector'("00000000000000000000000000000010"), A_WE_StdLogicVector((std_logic'((internal_pcp_cpu_instruction_master_granted_cfi_flash_0_s1)) = '1'), std_logic_vector'("00000000000000000000000000000010"), A_WE_StdLogicVector((std_logic'((internal_pcp_cpu_data_master_granted_DBC3C40_SRAM_0_avalon_tristate_slave)) = '1'), std_logic_vector'("00000000000000000000000000000010"), A_WE_StdLogicVector((std_logic'((internal_pcp_cpu_instruction_master_granted_DBC3C40_SRAM_0_avalon_tristate_slave)) = '1'), std_logic_vector'("00000000000000000000000000000010"), A_WE_StdLogicVector((std_logic'((internal_pcp_cpu_data_master_granted_cfi_flash_0_s1)) = '1'), std_logic_vector'("00000000000000000000000000000010"), A_WE_StdLogicVector((std_logic'((internal_pcp_cpu_instruction_master_granted_cfi_flash_0_s1)) = '1'), std_logic_vector'("00000000000000000000000000000010"), std_logic_vector'("00000000000000000000000000000001"))))))))), 2);
  --tri_state_bridge_0_avalon_slave_non_bursting_master_requests mux, which is an e_mux
  tri_state_bridge_0_avalon_slave_non_bursting_master_requests <= ((((((internal_pcp_cpu_data_master_requests_DBC3C40_SRAM_0_avalon_tristate_slave OR internal_pcp_cpu_instruction_master_requests_DBC3C40_SRAM_0_avalon_tristate_slave) OR internal_pcp_cpu_data_master_requests_cfi_flash_0_s1) OR internal_pcp_cpu_instruction_master_requests_cfi_flash_0_s1) OR internal_pcp_cpu_data_master_requests_DBC3C40_SRAM_0_avalon_tristate_slave) OR internal_pcp_cpu_instruction_master_requests_DBC3C40_SRAM_0_avalon_tristate_slave) OR internal_pcp_cpu_data_master_requests_cfi_flash_0_s1) OR internal_pcp_cpu_instruction_master_requests_cfi_flash_0_s1;
  --tri_state_bridge_0_avalon_slave_any_bursting_master_saved_grant mux, which is an e_mux
  tri_state_bridge_0_avalon_slave_any_bursting_master_saved_grant <= std_logic'('0');
  --tri_state_bridge_0_avalon_slave_arb_share_counter_next_value assignment, which is an e_assign
  tri_state_bridge_0_avalon_slave_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(tri_state_bridge_0_avalon_slave_firsttransfer) = '1'), (((std_logic_vector'("0000000000000000000000000000000") & (tri_state_bridge_0_avalon_slave_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(tri_state_bridge_0_avalon_slave_arb_share_counter)) = '1'), (((std_logic_vector'("0000000000000000000000000000000") & (tri_state_bridge_0_avalon_slave_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 2);
  --tri_state_bridge_0_avalon_slave_allgrants all slave grants, which is an e_mux
  tri_state_bridge_0_avalon_slave_allgrants <= (((((((or_reduce(tri_state_bridge_0_avalon_slave_grant_vector)) OR (or_reduce(tri_state_bridge_0_avalon_slave_grant_vector))) OR (or_reduce(tri_state_bridge_0_avalon_slave_grant_vector))) OR (or_reduce(tri_state_bridge_0_avalon_slave_grant_vector))) OR (or_reduce(tri_state_bridge_0_avalon_slave_grant_vector))) OR (or_reduce(tri_state_bridge_0_avalon_slave_grant_vector))) OR (or_reduce(tri_state_bridge_0_avalon_slave_grant_vector))) OR (or_reduce(tri_state_bridge_0_avalon_slave_grant_vector));
  --tri_state_bridge_0_avalon_slave_end_xfer assignment, which is an e_assign
  tri_state_bridge_0_avalon_slave_end_xfer <= NOT ((((DBC3C40_SRAM_0_avalon_tristate_slave_waits_for_read OR DBC3C40_SRAM_0_avalon_tristate_slave_waits_for_write) OR cfi_flash_0_s1_waits_for_read) OR cfi_flash_0_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_tri_state_bridge_0_avalon_slave arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_tri_state_bridge_0_avalon_slave <= tri_state_bridge_0_avalon_slave_end_xfer AND (((NOT tri_state_bridge_0_avalon_slave_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --tri_state_bridge_0_avalon_slave_arb_share_counter arbitration counter enable, which is an e_assign
  tri_state_bridge_0_avalon_slave_arb_counter_enable <= ((end_xfer_arb_share_counter_term_tri_state_bridge_0_avalon_slave AND tri_state_bridge_0_avalon_slave_allgrants)) OR ((end_xfer_arb_share_counter_term_tri_state_bridge_0_avalon_slave AND NOT tri_state_bridge_0_avalon_slave_non_bursting_master_requests));
  --tri_state_bridge_0_avalon_slave_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      tri_state_bridge_0_avalon_slave_arb_share_counter <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      if std_logic'(tri_state_bridge_0_avalon_slave_arb_counter_enable) = '1' then 
        tri_state_bridge_0_avalon_slave_arb_share_counter <= tri_state_bridge_0_avalon_slave_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --tri_state_bridge_0_avalon_slave_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      tri_state_bridge_0_avalon_slave_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((or_reduce(tri_state_bridge_0_avalon_slave_master_qreq_vector) AND end_xfer_arb_share_counter_term_tri_state_bridge_0_avalon_slave)) OR ((end_xfer_arb_share_counter_term_tri_state_bridge_0_avalon_slave AND NOT tri_state_bridge_0_avalon_slave_non_bursting_master_requests)))) = '1' then 
        tri_state_bridge_0_avalon_slave_slavearbiterlockenable <= or_reduce(tri_state_bridge_0_avalon_slave_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --pcp_cpu/data_master tri_state_bridge_0/avalon_slave arbiterlock, which is an e_assign
  pcp_cpu_data_master_arbiterlock <= tri_state_bridge_0_avalon_slave_slavearbiterlockenable AND pcp_cpu_data_master_continuerequest;
  --tri_state_bridge_0_avalon_slave_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  tri_state_bridge_0_avalon_slave_slavearbiterlockenable2 <= or_reduce(tri_state_bridge_0_avalon_slave_arb_share_counter_next_value);
  --pcp_cpu/data_master tri_state_bridge_0/avalon_slave arbiterlock2, which is an e_assign
  pcp_cpu_data_master_arbiterlock2 <= tri_state_bridge_0_avalon_slave_slavearbiterlockenable2 AND pcp_cpu_data_master_continuerequest;
  --pcp_cpu/instruction_master tri_state_bridge_0/avalon_slave arbiterlock, which is an e_assign
  pcp_cpu_instruction_master_arbiterlock <= tri_state_bridge_0_avalon_slave_slavearbiterlockenable AND pcp_cpu_instruction_master_continuerequest;
  --pcp_cpu/instruction_master tri_state_bridge_0/avalon_slave arbiterlock2, which is an e_assign
  pcp_cpu_instruction_master_arbiterlock2 <= tri_state_bridge_0_avalon_slave_slavearbiterlockenable2 AND pcp_cpu_instruction_master_continuerequest;
  --pcp_cpu/instruction_master granted DBC3C40_SRAM_0/avalon_tristate_slave last time, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      last_cycle_pcp_cpu_instruction_master_granted_slave_DBC3C40_SRAM_0_avalon_tristate_slave <= std_logic'('0');
    elsif clk'event and clk = '1' then
      last_cycle_pcp_cpu_instruction_master_granted_slave_DBC3C40_SRAM_0_avalon_tristate_slave <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(pcp_cpu_instruction_master_saved_grant_DBC3C40_SRAM_0_avalon_tristate_slave) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((tri_state_bridge_0_avalon_slave_arbitration_holdoff_internal OR NOT internal_pcp_cpu_instruction_master_requests_DBC3C40_SRAM_0_avalon_tristate_slave))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_pcp_cpu_instruction_master_granted_slave_DBC3C40_SRAM_0_avalon_tristate_slave))))));
    end if;

  end process;

  --pcp_cpu_instruction_master_continuerequest continued request, which is an e_mux
  pcp_cpu_instruction_master_continuerequest <= ((last_cycle_pcp_cpu_instruction_master_granted_slave_DBC3C40_SRAM_0_avalon_tristate_slave AND internal_pcp_cpu_instruction_master_requests_DBC3C40_SRAM_0_avalon_tristate_slave)) OR ((last_cycle_pcp_cpu_instruction_master_granted_slave_cfi_flash_0_s1 AND internal_pcp_cpu_instruction_master_requests_cfi_flash_0_s1));
  --tri_state_bridge_0_avalon_slave_any_continuerequest at least one master continues requesting, which is an e_mux
  tri_state_bridge_0_avalon_slave_any_continuerequest <= ((pcp_cpu_instruction_master_continuerequest OR pcp_cpu_instruction_master_continuerequest) OR pcp_cpu_data_master_continuerequest) OR pcp_cpu_data_master_continuerequest;
  internal_pcp_cpu_data_master_qualified_request_DBC3C40_SRAM_0_avalon_tristate_slave <= internal_pcp_cpu_data_master_requests_DBC3C40_SRAM_0_avalon_tristate_slave AND NOT (((((pcp_cpu_data_master_read AND (((tri_state_bridge_0_avalon_slave_write_pending OR (tri_state_bridge_0_avalon_slave_read_pending)) OR (or_reduce(pcp_cpu_data_master_read_data_valid_DBC3C40_SRAM_0_avalon_tristate_slave_shift_register)))))) OR (((((tri_state_bridge_0_avalon_slave_read_pending OR pcp_cpu_data_master_no_byte_enables_and_last_term) OR NOT(or_reduce(internal_pcp_cpu_data_master_byteenable_DBC3C40_SRAM_0_avalon_tristate_slave)))) AND pcp_cpu_data_master_write))) OR pcp_cpu_instruction_master_arbiterlock));
  --pcp_cpu_data_master_read_data_valid_DBC3C40_SRAM_0_avalon_tristate_slave_shift_register_in mux for readlatency shift register, which is an e_mux
  pcp_cpu_data_master_read_data_valid_DBC3C40_SRAM_0_avalon_tristate_slave_shift_register_in <= ((internal_pcp_cpu_data_master_granted_DBC3C40_SRAM_0_avalon_tristate_slave AND pcp_cpu_data_master_read) AND NOT DBC3C40_SRAM_0_avalon_tristate_slave_waits_for_read) AND NOT (or_reduce(pcp_cpu_data_master_read_data_valid_DBC3C40_SRAM_0_avalon_tristate_slave_shift_register));
  --shift register p1 pcp_cpu_data_master_read_data_valid_DBC3C40_SRAM_0_avalon_tristate_slave_shift_register in if flush, otherwise shift left, which is an e_mux
  p1_pcp_cpu_data_master_read_data_valid_DBC3C40_SRAM_0_avalon_tristate_slave_shift_register <= A_EXT ((pcp_cpu_data_master_read_data_valid_DBC3C40_SRAM_0_avalon_tristate_slave_shift_register & A_ToStdLogicVector(pcp_cpu_data_master_read_data_valid_DBC3C40_SRAM_0_avalon_tristate_slave_shift_register_in)), 2);
  --pcp_cpu_data_master_read_data_valid_DBC3C40_SRAM_0_avalon_tristate_slave_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pcp_cpu_data_master_read_data_valid_DBC3C40_SRAM_0_avalon_tristate_slave_shift_register <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      pcp_cpu_data_master_read_data_valid_DBC3C40_SRAM_0_avalon_tristate_slave_shift_register <= p1_pcp_cpu_data_master_read_data_valid_DBC3C40_SRAM_0_avalon_tristate_slave_shift_register;
    end if;

  end process;

  --local readdatavalid pcp_cpu_data_master_read_data_valid_DBC3C40_SRAM_0_avalon_tristate_slave, which is an e_mux
  pcp_cpu_data_master_read_data_valid_DBC3C40_SRAM_0_avalon_tristate_slave <= pcp_cpu_data_master_read_data_valid_DBC3C40_SRAM_0_avalon_tristate_slave_shift_register(1);
  --tri_state_bridge_0_data register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      internal_incoming_tri_state_bridge_0_data <= std_logic_vector'("0000000000000000");
    elsif clk'event and clk = '1' then
      internal_incoming_tri_state_bridge_0_data <= tri_state_bridge_0_data;
    end if;

  end process;

  --DBC3C40_SRAM_0_avalon_tristate_slave_with_write_latency assignment, which is an e_assign
  DBC3C40_SRAM_0_avalon_tristate_slave_with_write_latency <= in_a_write_cycle AND ((internal_pcp_cpu_data_master_qualified_request_DBC3C40_SRAM_0_avalon_tristate_slave OR internal_pcp_cpu_instruction_master_qualified_request_DBC3C40_SRAM_0_avalon_tristate_slave));
  --time to write the data, which is an e_mux
  time_to_write <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((DBC3C40_SRAM_0_avalon_tristate_slave_with_write_latency)) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'((cfi_flash_0_s1_with_write_latency)) = '1'), std_logic_vector'("00000000000000000000000000000001"), std_logic_vector'("00000000000000000000000000000000"))));
  --d1_outgoing_tri_state_bridge_0_data register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_outgoing_tri_state_bridge_0_data <= std_logic_vector'("0000000000000000");
    elsif clk'event and clk = '1' then
      d1_outgoing_tri_state_bridge_0_data <= outgoing_tri_state_bridge_0_data;
    end if;

  end process;

  --write cycle delayed by 1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_in_a_write_cycle <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_in_a_write_cycle <= time_to_write;
    end if;

  end process;

  --d1_outgoing_tri_state_bridge_0_data tristate driver, which is an e_assign
  tri_state_bridge_0_data <= A_WE_StdLogicVector((std_logic'((d1_in_a_write_cycle)) = '1'), d1_outgoing_tri_state_bridge_0_data, A_REP(std_logic'('Z'), 16));
  --outgoing_tri_state_bridge_0_data mux, which is an e_mux
  outgoing_tri_state_bridge_0_data <= A_WE_StdLogicVector((std_logic'((internal_pcp_cpu_data_master_granted_DBC3C40_SRAM_0_avalon_tristate_slave)) = '1'), pcp_cpu_data_master_dbs_write_16, pcp_cpu_data_master_dbs_write_16);
  internal_pcp_cpu_data_master_requests_cfi_flash_0_s1 <= to_std_logic(((Std_Logic_Vector'(pcp_cpu_data_master_address_to_slave(25 DOWNTO 23) & std_logic_vector'("00000000000000000000000")) = std_logic_vector'("10000000000000000000000000")))) AND ((pcp_cpu_data_master_read OR pcp_cpu_data_master_write));
  --registered rdv signal_name registered_pcp_cpu_data_master_read_data_valid_cfi_flash_0_s1 assignment, which is an e_assign
  registered_pcp_cpu_data_master_read_data_valid_cfi_flash_0_s1 <= pcp_cpu_data_master_read_data_valid_cfi_flash_0_s1_shift_register(0);
  --pcp_cpu/instruction_master granted cfi_flash_0/s1 last time, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      last_cycle_pcp_cpu_instruction_master_granted_slave_cfi_flash_0_s1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      last_cycle_pcp_cpu_instruction_master_granted_slave_cfi_flash_0_s1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(pcp_cpu_instruction_master_saved_grant_cfi_flash_0_s1) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((tri_state_bridge_0_avalon_slave_arbitration_holdoff_internal OR NOT internal_pcp_cpu_instruction_master_requests_cfi_flash_0_s1))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_pcp_cpu_instruction_master_granted_slave_cfi_flash_0_s1))))));
    end if;

  end process;

  internal_pcp_cpu_data_master_qualified_request_cfi_flash_0_s1 <= internal_pcp_cpu_data_master_requests_cfi_flash_0_s1 AND NOT (((((pcp_cpu_data_master_read AND (((tri_state_bridge_0_avalon_slave_write_pending OR (tri_state_bridge_0_avalon_slave_read_pending)) OR (or_reduce(pcp_cpu_data_master_read_data_valid_cfi_flash_0_s1_shift_register)))))) OR (((((tri_state_bridge_0_avalon_slave_read_pending OR pcp_cpu_data_master_no_byte_enables_and_last_term) OR NOT(or_reduce(internal_pcp_cpu_data_master_byteenable_cfi_flash_0_s1)))) AND pcp_cpu_data_master_write))) OR pcp_cpu_instruction_master_arbiterlock));
  --pcp_cpu_data_master_read_data_valid_cfi_flash_0_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  pcp_cpu_data_master_read_data_valid_cfi_flash_0_s1_shift_register_in <= ((internal_pcp_cpu_data_master_granted_cfi_flash_0_s1 AND pcp_cpu_data_master_read) AND NOT cfi_flash_0_s1_waits_for_read) AND NOT (or_reduce(pcp_cpu_data_master_read_data_valid_cfi_flash_0_s1_shift_register));
  --shift register p1 pcp_cpu_data_master_read_data_valid_cfi_flash_0_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  p1_pcp_cpu_data_master_read_data_valid_cfi_flash_0_s1_shift_register <= A_EXT ((pcp_cpu_data_master_read_data_valid_cfi_flash_0_s1_shift_register & A_ToStdLogicVector(pcp_cpu_data_master_read_data_valid_cfi_flash_0_s1_shift_register_in)), 2);
  --pcp_cpu_data_master_read_data_valid_cfi_flash_0_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pcp_cpu_data_master_read_data_valid_cfi_flash_0_s1_shift_register <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      pcp_cpu_data_master_read_data_valid_cfi_flash_0_s1_shift_register <= p1_pcp_cpu_data_master_read_data_valid_cfi_flash_0_s1_shift_register;
    end if;

  end process;

  --local readdatavalid pcp_cpu_data_master_read_data_valid_cfi_flash_0_s1, which is an e_mux
  pcp_cpu_data_master_read_data_valid_cfi_flash_0_s1 <= pcp_cpu_data_master_read_data_valid_cfi_flash_0_s1_shift_register(1);
  --cfi_flash_0_s1_with_write_latency assignment, which is an e_assign
  cfi_flash_0_s1_with_write_latency <= in_a_write_cycle AND ((internal_pcp_cpu_data_master_qualified_request_cfi_flash_0_s1 OR internal_pcp_cpu_instruction_master_qualified_request_cfi_flash_0_s1));
  internal_pcp_cpu_instruction_master_requests_DBC3C40_SRAM_0_avalon_tristate_slave <= ((to_std_logic(((Std_Logic_Vector'(pcp_cpu_instruction_master_address_to_slave(25 DOWNTO 20) & std_logic_vector'("00000000000000000000")) = std_logic_vector'("00001000000000000000000000")))) AND (pcp_cpu_instruction_master_read))) AND pcp_cpu_instruction_master_read;
  --pcp_cpu/data_master granted DBC3C40_SRAM_0/avalon_tristate_slave last time, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      last_cycle_pcp_cpu_data_master_granted_slave_DBC3C40_SRAM_0_avalon_tristate_slave <= std_logic'('0');
    elsif clk'event and clk = '1' then
      last_cycle_pcp_cpu_data_master_granted_slave_DBC3C40_SRAM_0_avalon_tristate_slave <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(pcp_cpu_data_master_saved_grant_DBC3C40_SRAM_0_avalon_tristate_slave) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((tri_state_bridge_0_avalon_slave_arbitration_holdoff_internal OR NOT internal_pcp_cpu_data_master_requests_DBC3C40_SRAM_0_avalon_tristate_slave))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_pcp_cpu_data_master_granted_slave_DBC3C40_SRAM_0_avalon_tristate_slave))))));
    end if;

  end process;

  --pcp_cpu_data_master_continuerequest continued request, which is an e_mux
  pcp_cpu_data_master_continuerequest <= ((last_cycle_pcp_cpu_data_master_granted_slave_DBC3C40_SRAM_0_avalon_tristate_slave AND internal_pcp_cpu_data_master_requests_DBC3C40_SRAM_0_avalon_tristate_slave)) OR ((last_cycle_pcp_cpu_data_master_granted_slave_cfi_flash_0_s1 AND internal_pcp_cpu_data_master_requests_cfi_flash_0_s1));
  internal_pcp_cpu_instruction_master_qualified_request_DBC3C40_SRAM_0_avalon_tristate_slave <= internal_pcp_cpu_instruction_master_requests_DBC3C40_SRAM_0_avalon_tristate_slave AND NOT ((((pcp_cpu_instruction_master_read AND (((tri_state_bridge_0_avalon_slave_write_pending OR (tri_state_bridge_0_avalon_slave_read_pending)) OR to_std_logic(((std_logic_vector'("00000000000000000000000000000010")<(std_logic_vector'("000000000000000000000000000000") & (pcp_cpu_instruction_master_latency_counter))))))))) OR pcp_cpu_data_master_arbiterlock));
  --pcp_cpu_instruction_master_read_data_valid_DBC3C40_SRAM_0_avalon_tristate_slave_shift_register_in mux for readlatency shift register, which is an e_mux
  pcp_cpu_instruction_master_read_data_valid_DBC3C40_SRAM_0_avalon_tristate_slave_shift_register_in <= (internal_pcp_cpu_instruction_master_granted_DBC3C40_SRAM_0_avalon_tristate_slave AND pcp_cpu_instruction_master_read) AND NOT DBC3C40_SRAM_0_avalon_tristate_slave_waits_for_read;
  --shift register p1 pcp_cpu_instruction_master_read_data_valid_DBC3C40_SRAM_0_avalon_tristate_slave_shift_register in if flush, otherwise shift left, which is an e_mux
  p1_pcp_cpu_instruction_master_read_data_valid_DBC3C40_SRAM_0_avalon_tristate_slave_shift_register <= A_EXT ((pcp_cpu_instruction_master_read_data_valid_DBC3C40_SRAM_0_avalon_tristate_slave_shift_register & A_ToStdLogicVector(pcp_cpu_instruction_master_read_data_valid_DBC3C40_SRAM_0_avalon_tristate_slave_shift_register_in)), 2);
  --pcp_cpu_instruction_master_read_data_valid_DBC3C40_SRAM_0_avalon_tristate_slave_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pcp_cpu_instruction_master_read_data_valid_DBC3C40_SRAM_0_avalon_tristate_slave_shift_register <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      pcp_cpu_instruction_master_read_data_valid_DBC3C40_SRAM_0_avalon_tristate_slave_shift_register <= p1_pcp_cpu_instruction_master_read_data_valid_DBC3C40_SRAM_0_avalon_tristate_slave_shift_register;
    end if;

  end process;

  --local readdatavalid pcp_cpu_instruction_master_read_data_valid_DBC3C40_SRAM_0_avalon_tristate_slave, which is an e_mux
  pcp_cpu_instruction_master_read_data_valid_DBC3C40_SRAM_0_avalon_tristate_slave <= pcp_cpu_instruction_master_read_data_valid_DBC3C40_SRAM_0_avalon_tristate_slave_shift_register(1);
  internal_pcp_cpu_instruction_master_requests_cfi_flash_0_s1 <= ((to_std_logic(((Std_Logic_Vector'(pcp_cpu_instruction_master_address_to_slave(25 DOWNTO 23) & std_logic_vector'("00000000000000000000000")) = std_logic_vector'("10000000000000000000000000")))) AND (pcp_cpu_instruction_master_read))) AND pcp_cpu_instruction_master_read;
  --pcp_cpu/data_master granted cfi_flash_0/s1 last time, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      last_cycle_pcp_cpu_data_master_granted_slave_cfi_flash_0_s1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      last_cycle_pcp_cpu_data_master_granted_slave_cfi_flash_0_s1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(pcp_cpu_data_master_saved_grant_cfi_flash_0_s1) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((tri_state_bridge_0_avalon_slave_arbitration_holdoff_internal OR NOT internal_pcp_cpu_data_master_requests_cfi_flash_0_s1))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_pcp_cpu_data_master_granted_slave_cfi_flash_0_s1))))));
    end if;

  end process;

  internal_pcp_cpu_instruction_master_qualified_request_cfi_flash_0_s1 <= internal_pcp_cpu_instruction_master_requests_cfi_flash_0_s1 AND NOT ((((pcp_cpu_instruction_master_read AND (((tri_state_bridge_0_avalon_slave_write_pending OR (tri_state_bridge_0_avalon_slave_read_pending)) OR to_std_logic(((std_logic_vector'("00000000000000000000000000000010")<(std_logic_vector'("000000000000000000000000000000") & (pcp_cpu_instruction_master_latency_counter))))))))) OR pcp_cpu_data_master_arbiterlock));
  --pcp_cpu_instruction_master_read_data_valid_cfi_flash_0_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  pcp_cpu_instruction_master_read_data_valid_cfi_flash_0_s1_shift_register_in <= (internal_pcp_cpu_instruction_master_granted_cfi_flash_0_s1 AND pcp_cpu_instruction_master_read) AND NOT cfi_flash_0_s1_waits_for_read;
  --shift register p1 pcp_cpu_instruction_master_read_data_valid_cfi_flash_0_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  p1_pcp_cpu_instruction_master_read_data_valid_cfi_flash_0_s1_shift_register <= A_EXT ((pcp_cpu_instruction_master_read_data_valid_cfi_flash_0_s1_shift_register & A_ToStdLogicVector(pcp_cpu_instruction_master_read_data_valid_cfi_flash_0_s1_shift_register_in)), 2);
  --pcp_cpu_instruction_master_read_data_valid_cfi_flash_0_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pcp_cpu_instruction_master_read_data_valid_cfi_flash_0_s1_shift_register <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      pcp_cpu_instruction_master_read_data_valid_cfi_flash_0_s1_shift_register <= p1_pcp_cpu_instruction_master_read_data_valid_cfi_flash_0_s1_shift_register;
    end if;

  end process;

  --local readdatavalid pcp_cpu_instruction_master_read_data_valid_cfi_flash_0_s1, which is an e_mux
  pcp_cpu_instruction_master_read_data_valid_cfi_flash_0_s1 <= pcp_cpu_instruction_master_read_data_valid_cfi_flash_0_s1_shift_register(1);
  --allow new arb cycle for tri_state_bridge_0/avalon_slave, which is an e_assign
  tri_state_bridge_0_avalon_slave_allow_new_arb_cycle <= NOT pcp_cpu_data_master_arbiterlock AND NOT pcp_cpu_instruction_master_arbiterlock;
  --pcp_cpu/instruction_master assignment into master qualified-requests vector for DBC3C40_SRAM_0/avalon_tristate_slave, which is an e_assign
  tri_state_bridge_0_avalon_slave_master_qreq_vector(0) <= internal_pcp_cpu_instruction_master_qualified_request_DBC3C40_SRAM_0_avalon_tristate_slave;
  --pcp_cpu/instruction_master grant DBC3C40_SRAM_0/avalon_tristate_slave, which is an e_assign
  internal_pcp_cpu_instruction_master_granted_DBC3C40_SRAM_0_avalon_tristate_slave <= tri_state_bridge_0_avalon_slave_grant_vector(0);
  --pcp_cpu/instruction_master saved-grant DBC3C40_SRAM_0/avalon_tristate_slave, which is an e_assign
  pcp_cpu_instruction_master_saved_grant_DBC3C40_SRAM_0_avalon_tristate_slave <= tri_state_bridge_0_avalon_slave_arb_winner(0) AND internal_pcp_cpu_instruction_master_requests_DBC3C40_SRAM_0_avalon_tristate_slave;
  --pcp_cpu/data_master assignment into master qualified-requests vector for DBC3C40_SRAM_0/avalon_tristate_slave, which is an e_assign
  tri_state_bridge_0_avalon_slave_master_qreq_vector(1) <= internal_pcp_cpu_data_master_qualified_request_DBC3C40_SRAM_0_avalon_tristate_slave;
  --pcp_cpu/data_master grant DBC3C40_SRAM_0/avalon_tristate_slave, which is an e_assign
  internal_pcp_cpu_data_master_granted_DBC3C40_SRAM_0_avalon_tristate_slave <= tri_state_bridge_0_avalon_slave_grant_vector(1);
  --pcp_cpu/data_master saved-grant DBC3C40_SRAM_0/avalon_tristate_slave, which is an e_assign
  pcp_cpu_data_master_saved_grant_DBC3C40_SRAM_0_avalon_tristate_slave <= tri_state_bridge_0_avalon_slave_arb_winner(1) AND internal_pcp_cpu_data_master_requests_DBC3C40_SRAM_0_avalon_tristate_slave;
  --pcp_cpu/instruction_master assignment into master qualified-requests vector for cfi_flash_0/s1, which is an e_assign
  tri_state_bridge_0_avalon_slave_master_qreq_vector(2) <= internal_pcp_cpu_instruction_master_qualified_request_cfi_flash_0_s1;
  --pcp_cpu/instruction_master grant cfi_flash_0/s1, which is an e_assign
  internal_pcp_cpu_instruction_master_granted_cfi_flash_0_s1 <= tri_state_bridge_0_avalon_slave_grant_vector(2);
  --pcp_cpu/instruction_master saved-grant cfi_flash_0/s1, which is an e_assign
  pcp_cpu_instruction_master_saved_grant_cfi_flash_0_s1 <= tri_state_bridge_0_avalon_slave_arb_winner(2) AND internal_pcp_cpu_instruction_master_requests_cfi_flash_0_s1;
  --pcp_cpu/data_master assignment into master qualified-requests vector for cfi_flash_0/s1, which is an e_assign
  tri_state_bridge_0_avalon_slave_master_qreq_vector(3) <= internal_pcp_cpu_data_master_qualified_request_cfi_flash_0_s1;
  --pcp_cpu/data_master grant cfi_flash_0/s1, which is an e_assign
  internal_pcp_cpu_data_master_granted_cfi_flash_0_s1 <= tri_state_bridge_0_avalon_slave_grant_vector(3);
  --pcp_cpu/data_master saved-grant cfi_flash_0/s1, which is an e_assign
  pcp_cpu_data_master_saved_grant_cfi_flash_0_s1 <= tri_state_bridge_0_avalon_slave_arb_winner(3) AND internal_pcp_cpu_data_master_requests_cfi_flash_0_s1;
  --tri_state_bridge_0/avalon_slave chosen-master double-vector, which is an e_assign
  tri_state_bridge_0_avalon_slave_chosen_master_double_vector <= A_EXT (((std_logic_vector'("0") & ((tri_state_bridge_0_avalon_slave_master_qreq_vector & tri_state_bridge_0_avalon_slave_master_qreq_vector))) AND (((std_logic_vector'("0") & (Std_Logic_Vector'(NOT tri_state_bridge_0_avalon_slave_master_qreq_vector & NOT tri_state_bridge_0_avalon_slave_master_qreq_vector))) + (std_logic_vector'("00000") & (tri_state_bridge_0_avalon_slave_arb_addend))))), 8);
  --stable onehot encoding of arb winner
  tri_state_bridge_0_avalon_slave_arb_winner <= A_WE_StdLogicVector((std_logic'(((tri_state_bridge_0_avalon_slave_allow_new_arb_cycle AND or_reduce(tri_state_bridge_0_avalon_slave_grant_vector)))) = '1'), tri_state_bridge_0_avalon_slave_grant_vector, tri_state_bridge_0_avalon_slave_saved_chosen_master_vector);
  --saved tri_state_bridge_0_avalon_slave_grant_vector, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      tri_state_bridge_0_avalon_slave_saved_chosen_master_vector <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'(tri_state_bridge_0_avalon_slave_allow_new_arb_cycle) = '1' then 
        tri_state_bridge_0_avalon_slave_saved_chosen_master_vector <= A_WE_StdLogicVector((std_logic'(or_reduce(tri_state_bridge_0_avalon_slave_grant_vector)) = '1'), tri_state_bridge_0_avalon_slave_grant_vector, tri_state_bridge_0_avalon_slave_saved_chosen_master_vector);
      end if;
    end if;

  end process;

  --onehot encoding of chosen master
  tri_state_bridge_0_avalon_slave_grant_vector <= Std_Logic_Vector'(A_ToStdLogicVector(((tri_state_bridge_0_avalon_slave_chosen_master_double_vector(3) OR tri_state_bridge_0_avalon_slave_chosen_master_double_vector(7)))) & A_ToStdLogicVector(((tri_state_bridge_0_avalon_slave_chosen_master_double_vector(2) OR tri_state_bridge_0_avalon_slave_chosen_master_double_vector(6)))) & A_ToStdLogicVector(((tri_state_bridge_0_avalon_slave_chosen_master_double_vector(1) OR tri_state_bridge_0_avalon_slave_chosen_master_double_vector(5)))) & A_ToStdLogicVector(((tri_state_bridge_0_avalon_slave_chosen_master_double_vector(0) OR tri_state_bridge_0_avalon_slave_chosen_master_double_vector(4)))));
  --tri_state_bridge_0/avalon_slave chosen master rotated left, which is an e_assign
  tri_state_bridge_0_avalon_slave_chosen_master_rot_left <= A_EXT (A_WE_StdLogicVector((((A_SLL(tri_state_bridge_0_avalon_slave_arb_winner,std_logic_vector'("00000000000000000000000000000001")))) /= std_logic_vector'("0000")), (std_logic_vector'("0000000000000000000000000000") & ((A_SLL(tri_state_bridge_0_avalon_slave_arb_winner,std_logic_vector'("00000000000000000000000000000001"))))), std_logic_vector'("00000000000000000000000000000001")), 4);
  --tri_state_bridge_0/avalon_slave's addend for next-master-grant
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      tri_state_bridge_0_avalon_slave_arb_addend <= std_logic_vector'("0001");
    elsif clk'event and clk = '1' then
      if std_logic'(or_reduce(tri_state_bridge_0_avalon_slave_grant_vector)) = '1' then 
        tri_state_bridge_0_avalon_slave_arb_addend <= A_WE_StdLogicVector((std_logic'(tri_state_bridge_0_avalon_slave_end_xfer) = '1'), tri_state_bridge_0_avalon_slave_chosen_master_rot_left, tri_state_bridge_0_avalon_slave_grant_vector);
      end if;
    end if;

  end process;

  p1_ncs_to_the_DBC3C40_SRAM_0 <= NOT ((internal_pcp_cpu_data_master_granted_DBC3C40_SRAM_0_avalon_tristate_slave OR internal_pcp_cpu_instruction_master_granted_DBC3C40_SRAM_0_avalon_tristate_slave));
  --tri_state_bridge_0_avalon_slave_firsttransfer first transaction, which is an e_assign
  tri_state_bridge_0_avalon_slave_firsttransfer <= A_WE_StdLogic((std_logic'(tri_state_bridge_0_avalon_slave_begins_xfer) = '1'), tri_state_bridge_0_avalon_slave_unreg_firsttransfer, tri_state_bridge_0_avalon_slave_reg_firsttransfer);
  --tri_state_bridge_0_avalon_slave_unreg_firsttransfer first transaction, which is an e_assign
  tri_state_bridge_0_avalon_slave_unreg_firsttransfer <= NOT ((tri_state_bridge_0_avalon_slave_slavearbiterlockenable AND tri_state_bridge_0_avalon_slave_any_continuerequest));
  --tri_state_bridge_0_avalon_slave_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      tri_state_bridge_0_avalon_slave_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(tri_state_bridge_0_avalon_slave_begins_xfer) = '1' then 
        tri_state_bridge_0_avalon_slave_reg_firsttransfer <= tri_state_bridge_0_avalon_slave_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --tri_state_bridge_0_avalon_slave_beginbursttransfer_internal begin burst transfer, which is an e_assign
  tri_state_bridge_0_avalon_slave_beginbursttransfer_internal <= tri_state_bridge_0_avalon_slave_begins_xfer;
  --tri_state_bridge_0_avalon_slave_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  tri_state_bridge_0_avalon_slave_arbitration_holdoff_internal <= tri_state_bridge_0_avalon_slave_begins_xfer AND tri_state_bridge_0_avalon_slave_firsttransfer;
  --~tri_state_bridge_0_readn of type read to ~p1_tri_state_bridge_0_readn, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      tri_state_bridge_0_readn <= Vector_To_Std_Logic(NOT std_logic_vector'("00000000000000000000000000000000"));
    elsif clk'event and clk = '1' then
      tri_state_bridge_0_readn <= p1_tri_state_bridge_0_readn;
    end if;

  end process;

  --~p1_tri_state_bridge_0_readn assignment, which is an e_mux
  p1_tri_state_bridge_0_readn <= NOT ((((((internal_pcp_cpu_data_master_granted_DBC3C40_SRAM_0_avalon_tristate_slave AND pcp_cpu_data_master_read)) OR ((internal_pcp_cpu_instruction_master_granted_DBC3C40_SRAM_0_avalon_tristate_slave AND pcp_cpu_instruction_master_read)))) OR ((((((internal_pcp_cpu_data_master_granted_cfi_flash_0_s1 AND pcp_cpu_data_master_read)) OR ((internal_pcp_cpu_instruction_master_granted_cfi_flash_0_s1 AND pcp_cpu_instruction_master_read)))) AND NOT tri_state_bridge_0_avalon_slave_begins_xfer))));
  --~tri_state_bridge_0_writen of type write to ~p1_tri_state_bridge_0_writen, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      tri_state_bridge_0_writen <= Vector_To_Std_Logic(NOT std_logic_vector'("00000000000000000000000000000000"));
    elsif clk'event and clk = '1' then
      tri_state_bridge_0_writen <= p1_tri_state_bridge_0_writen;
    end if;

  end process;

  --~ben_to_the_DBC3C40_SRAM_0 of type byteenable to ~p1_ben_to_the_DBC3C40_SRAM_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      ben_to_the_DBC3C40_SRAM_0 <= A_EXT (NOT std_logic_vector'("00000000000000000000000000000000"), 2);
    elsif clk'event and clk = '1' then
      ben_to_the_DBC3C40_SRAM_0 <= p1_ben_to_the_DBC3C40_SRAM_0;
    end if;

  end process;

  --~p1_tri_state_bridge_0_writen assignment, which is an e_mux
  p1_tri_state_bridge_0_writen <= NOT ((((((internal_pcp_cpu_data_master_granted_DBC3C40_SRAM_0_avalon_tristate_slave AND pcp_cpu_data_master_write)) AND ((tri_state_bridge_0_avalon_slave_begins_xfer OR to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(DBC3C40_SRAM_0_avalon_tristate_slave_wait_counter)))>=std_logic_vector'("00000000000000000000000000000001")))))))) OR (((((internal_pcp_cpu_data_master_granted_cfi_flash_0_s1 AND pcp_cpu_data_master_write)) AND NOT tri_state_bridge_0_avalon_slave_begins_xfer) AND to_std_logic((((std_logic_vector'("0000000000000000000000000000") & (cfi_flash_0_s1_wait_counter))>=std_logic_vector'("00000000000000000000000000000001"))))))));
  --tri_state_bridge_0_address of type address to p1_tri_state_bridge_0_address, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      tri_state_bridge_0_address <= std_logic_vector'("00000000000000000000000");
    elsif clk'event and clk = '1' then
      tri_state_bridge_0_address <= p1_tri_state_bridge_0_address;
    end if;

  end process;

  --p1_tri_state_bridge_0_address mux, which is an e_mux
  p1_tri_state_bridge_0_address <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_pcp_cpu_data_master_granted_DBC3C40_SRAM_0_avalon_tristate_slave)) = '1'), (Std_Logic_Vector'(A_SRL(pcp_cpu_data_master_address_to_slave,std_logic_vector'("00000000000000000000000000000010")) & A_ToStdLogicVector(pcp_cpu_data_master_dbs_address(1)) & A_ToStdLogicVector(std_logic'('0')))), A_WE_StdLogicVector((std_logic'((internal_pcp_cpu_instruction_master_granted_DBC3C40_SRAM_0_avalon_tristate_slave)) = '1'), (Std_Logic_Vector'(A_SRL(pcp_cpu_instruction_master_address_to_slave,std_logic_vector'("00000000000000000000000000000010")) & A_ToStdLogicVector(pcp_cpu_instruction_master_dbs_address(1)) & A_ToStdLogicVector(std_logic'('0')))), A_WE_StdLogicVector((std_logic'((internal_pcp_cpu_data_master_granted_cfi_flash_0_s1)) = '1'), (Std_Logic_Vector'(A_SRL(pcp_cpu_data_master_address_to_slave,std_logic_vector'("00000000000000000000000000000010")) & A_ToStdLogicVector(pcp_cpu_data_master_dbs_address(1)) & A_ToStdLogicVector(std_logic'('0')))), (Std_Logic_Vector'(A_SRL(pcp_cpu_instruction_master_address_to_slave,std_logic_vector'("00000000000000000000000000000010")) & A_ToStdLogicVector(pcp_cpu_instruction_master_dbs_address(1)) & A_ToStdLogicVector(std_logic'('0'))))))), 23);
  --d1_tri_state_bridge_0_avalon_slave_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_tri_state_bridge_0_avalon_slave_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_tri_state_bridge_0_avalon_slave_end_xfer <= tri_state_bridge_0_avalon_slave_end_xfer;
    end if;

  end process;

  --DBC3C40_SRAM_0_avalon_tristate_slave_waits_for_read in a cycle, which is an e_mux
  DBC3C40_SRAM_0_avalon_tristate_slave_waits_for_read <= DBC3C40_SRAM_0_avalon_tristate_slave_in_a_read_cycle AND wait_for_DBC3C40_SRAM_0_avalon_tristate_slave_counter;
  --DBC3C40_SRAM_0_avalon_tristate_slave_in_a_read_cycle assignment, which is an e_assign
  DBC3C40_SRAM_0_avalon_tristate_slave_in_a_read_cycle <= ((internal_pcp_cpu_data_master_granted_DBC3C40_SRAM_0_avalon_tristate_slave AND pcp_cpu_data_master_read)) OR ((internal_pcp_cpu_instruction_master_granted_DBC3C40_SRAM_0_avalon_tristate_slave AND pcp_cpu_instruction_master_read));
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= DBC3C40_SRAM_0_avalon_tristate_slave_in_a_read_cycle OR cfi_flash_0_s1_in_a_read_cycle;
  --DBC3C40_SRAM_0_avalon_tristate_slave_waits_for_write in a cycle, which is an e_mux
  DBC3C40_SRAM_0_avalon_tristate_slave_waits_for_write <= DBC3C40_SRAM_0_avalon_tristate_slave_in_a_write_cycle AND wait_for_DBC3C40_SRAM_0_avalon_tristate_slave_counter;
  --DBC3C40_SRAM_0_avalon_tristate_slave_in_a_write_cycle assignment, which is an e_assign
  DBC3C40_SRAM_0_avalon_tristate_slave_in_a_write_cycle <= internal_pcp_cpu_data_master_granted_DBC3C40_SRAM_0_avalon_tristate_slave AND pcp_cpu_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= DBC3C40_SRAM_0_avalon_tristate_slave_in_a_write_cycle OR cfi_flash_0_s1_in_a_write_cycle;
  internal_DBC3C40_SRAM_0_avalon_tristate_slave_wait_counter_eq_0 <= to_std_logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(DBC3C40_SRAM_0_avalon_tristate_slave_wait_counter))) = std_logic_vector'("00000000000000000000000000000000")));
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      DBC3C40_SRAM_0_avalon_tristate_slave_wait_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      DBC3C40_SRAM_0_avalon_tristate_slave_wait_counter <= DBC3C40_SRAM_0_avalon_tristate_slave_counter_load_value;
    end if;

  end process;

  DBC3C40_SRAM_0_avalon_tristate_slave_counter_load_value <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(((DBC3C40_SRAM_0_avalon_tristate_slave_in_a_write_cycle AND tri_state_bridge_0_avalon_slave_begins_xfer))) = '1'), std_logic_vector'("000000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((DBC3C40_SRAM_0_avalon_tristate_slave_in_a_read_cycle AND tri_state_bridge_0_avalon_slave_begins_xfer))) = '1'), std_logic_vector'("000000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'((NOT internal_DBC3C40_SRAM_0_avalon_tristate_slave_wait_counter_eq_0)) = '1'), ((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(DBC3C40_SRAM_0_avalon_tristate_slave_wait_counter))) - std_logic_vector'("000000000000000000000000000000001")), std_logic_vector'("000000000000000000000000000000000")))));
  wait_for_DBC3C40_SRAM_0_avalon_tristate_slave_counter <= tri_state_bridge_0_avalon_slave_begins_xfer OR NOT internal_DBC3C40_SRAM_0_avalon_tristate_slave_wait_counter_eq_0;
  --~p1_ben_to_the_DBC3C40_SRAM_0 byte enable port mux, which is an e_mux
  p1_ben_to_the_DBC3C40_SRAM_0 <= A_EXT (NOT (A_WE_StdLogicVector((std_logic'((internal_pcp_cpu_data_master_granted_DBC3C40_SRAM_0_avalon_tristate_slave)) = '1'), (std_logic_vector'("000000000000000000000000000000") & (internal_pcp_cpu_data_master_byteenable_DBC3C40_SRAM_0_avalon_tristate_slave)), -SIGNED(std_logic_vector'("00000000000000000000000000000001")))), 2);
  (pcp_cpu_data_master_byteenable_DBC3C40_SRAM_0_avalon_tristate_slave_segment_1(1), pcp_cpu_data_master_byteenable_DBC3C40_SRAM_0_avalon_tristate_slave_segment_1(0), pcp_cpu_data_master_byteenable_DBC3C40_SRAM_0_avalon_tristate_slave_segment_0(1), pcp_cpu_data_master_byteenable_DBC3C40_SRAM_0_avalon_tristate_slave_segment_0(0)) <= pcp_cpu_data_master_byteenable;
  internal_pcp_cpu_data_master_byteenable_DBC3C40_SRAM_0_avalon_tristate_slave <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pcp_cpu_data_master_dbs_address(1)))) = std_logic_vector'("00000000000000000000000000000000"))), pcp_cpu_data_master_byteenable_DBC3C40_SRAM_0_avalon_tristate_slave_segment_0, pcp_cpu_data_master_byteenable_DBC3C40_SRAM_0_avalon_tristate_slave_segment_1);
  p1_select_n_to_the_cfi_flash_0 <= NOT ((internal_pcp_cpu_data_master_granted_cfi_flash_0_s1 OR internal_pcp_cpu_instruction_master_granted_cfi_flash_0_s1));
  --cfi_flash_0_s1_wait_counter_eq_1 assignment, which is an e_assign
  cfi_flash_0_s1_wait_counter_eq_1 <= to_std_logic(((std_logic_vector'("0000000000000000000000000000") & (cfi_flash_0_s1_wait_counter)) = std_logic_vector'("00000000000000000000000000000001")));
  --cfi_flash_0_s1_waits_for_read in a cycle, which is an e_mux
  cfi_flash_0_s1_waits_for_read <= cfi_flash_0_s1_in_a_read_cycle AND wait_for_cfi_flash_0_s1_counter;
  --cfi_flash_0_s1_in_a_read_cycle assignment, which is an e_assign
  cfi_flash_0_s1_in_a_read_cycle <= ((internal_pcp_cpu_data_master_granted_cfi_flash_0_s1 AND pcp_cpu_data_master_read)) OR ((internal_pcp_cpu_instruction_master_granted_cfi_flash_0_s1 AND pcp_cpu_instruction_master_read));
  --cfi_flash_0_s1_waits_for_write in a cycle, which is an e_mux
  cfi_flash_0_s1_waits_for_write <= cfi_flash_0_s1_in_a_write_cycle AND wait_for_cfi_flash_0_s1_counter;
  --cfi_flash_0_s1_in_a_write_cycle assignment, which is an e_assign
  cfi_flash_0_s1_in_a_write_cycle <= internal_pcp_cpu_data_master_granted_cfi_flash_0_s1 AND pcp_cpu_data_master_write;
  internal_cfi_flash_0_s1_wait_counter_eq_0 <= to_std_logic(((std_logic_vector'("0000000000000000000000000000") & (cfi_flash_0_s1_wait_counter)) = std_logic_vector'("00000000000000000000000000000000")));
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      cfi_flash_0_s1_wait_counter <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      cfi_flash_0_s1_wait_counter <= cfi_flash_0_s1_counter_load_value;
    end if;

  end process;

  cfi_flash_0_s1_counter_load_value <= A_EXT (A_WE_StdLogicVector((std_logic'(((cfi_flash_0_s1_in_a_write_cycle AND tri_state_bridge_0_avalon_slave_begins_xfer))) = '1'), std_logic_vector'("000000000000000000000000000001001"), A_WE_StdLogicVector((std_logic'(((cfi_flash_0_s1_in_a_read_cycle AND tri_state_bridge_0_avalon_slave_begins_xfer))) = '1'), std_logic_vector'("000000000000000000000000000001000"), A_WE_StdLogicVector((std_logic'((NOT internal_cfi_flash_0_s1_wait_counter_eq_0)) = '1'), ((std_logic_vector'("00000000000000000000000000000") & (cfi_flash_0_s1_wait_counter)) - std_logic_vector'("000000000000000000000000000000001")), std_logic_vector'("000000000000000000000000000000000")))), 4);
  wait_for_cfi_flash_0_s1_counter <= tri_state_bridge_0_avalon_slave_begins_xfer OR NOT internal_cfi_flash_0_s1_wait_counter_eq_0;
  (pcp_cpu_data_master_byteenable_cfi_flash_0_s1_segment_1(1), pcp_cpu_data_master_byteenable_cfi_flash_0_s1_segment_1(0), pcp_cpu_data_master_byteenable_cfi_flash_0_s1_segment_0(1), pcp_cpu_data_master_byteenable_cfi_flash_0_s1_segment_0(0)) <= pcp_cpu_data_master_byteenable;
  internal_pcp_cpu_data_master_byteenable_cfi_flash_0_s1 <= A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pcp_cpu_data_master_dbs_address(1)))) = std_logic_vector'("00000000000000000000000000000000"))), pcp_cpu_data_master_byteenable_cfi_flash_0_s1_segment_0, pcp_cpu_data_master_byteenable_cfi_flash_0_s1_segment_1);
  --vhdl renameroo for output signals
  DBC3C40_SRAM_0_avalon_tristate_slave_wait_counter_eq_0 <= internal_DBC3C40_SRAM_0_avalon_tristate_slave_wait_counter_eq_0;
  --vhdl renameroo for output signals
  cfi_flash_0_s1_wait_counter_eq_0 <= internal_cfi_flash_0_s1_wait_counter_eq_0;
  --vhdl renameroo for output signals
  incoming_tri_state_bridge_0_data <= internal_incoming_tri_state_bridge_0_data;
  --vhdl renameroo for output signals
  pcp_cpu_data_master_byteenable_DBC3C40_SRAM_0_avalon_tristate_slave <= internal_pcp_cpu_data_master_byteenable_DBC3C40_SRAM_0_avalon_tristate_slave;
  --vhdl renameroo for output signals
  pcp_cpu_data_master_byteenable_cfi_flash_0_s1 <= internal_pcp_cpu_data_master_byteenable_cfi_flash_0_s1;
  --vhdl renameroo for output signals
  pcp_cpu_data_master_granted_DBC3C40_SRAM_0_avalon_tristate_slave <= internal_pcp_cpu_data_master_granted_DBC3C40_SRAM_0_avalon_tristate_slave;
  --vhdl renameroo for output signals
  pcp_cpu_data_master_granted_cfi_flash_0_s1 <= internal_pcp_cpu_data_master_granted_cfi_flash_0_s1;
  --vhdl renameroo for output signals
  pcp_cpu_data_master_qualified_request_DBC3C40_SRAM_0_avalon_tristate_slave <= internal_pcp_cpu_data_master_qualified_request_DBC3C40_SRAM_0_avalon_tristate_slave;
  --vhdl renameroo for output signals
  pcp_cpu_data_master_qualified_request_cfi_flash_0_s1 <= internal_pcp_cpu_data_master_qualified_request_cfi_flash_0_s1;
  --vhdl renameroo for output signals
  pcp_cpu_data_master_requests_DBC3C40_SRAM_0_avalon_tristate_slave <= internal_pcp_cpu_data_master_requests_DBC3C40_SRAM_0_avalon_tristate_slave;
  --vhdl renameroo for output signals
  pcp_cpu_data_master_requests_cfi_flash_0_s1 <= internal_pcp_cpu_data_master_requests_cfi_flash_0_s1;
  --vhdl renameroo for output signals
  pcp_cpu_instruction_master_granted_DBC3C40_SRAM_0_avalon_tristate_slave <= internal_pcp_cpu_instruction_master_granted_DBC3C40_SRAM_0_avalon_tristate_slave;
  --vhdl renameroo for output signals
  pcp_cpu_instruction_master_granted_cfi_flash_0_s1 <= internal_pcp_cpu_instruction_master_granted_cfi_flash_0_s1;
  --vhdl renameroo for output signals
  pcp_cpu_instruction_master_qualified_request_DBC3C40_SRAM_0_avalon_tristate_slave <= internal_pcp_cpu_instruction_master_qualified_request_DBC3C40_SRAM_0_avalon_tristate_slave;
  --vhdl renameroo for output signals
  pcp_cpu_instruction_master_qualified_request_cfi_flash_0_s1 <= internal_pcp_cpu_instruction_master_qualified_request_cfi_flash_0_s1;
  --vhdl renameroo for output signals
  pcp_cpu_instruction_master_requests_DBC3C40_SRAM_0_avalon_tristate_slave <= internal_pcp_cpu_instruction_master_requests_DBC3C40_SRAM_0_avalon_tristate_slave;
  --vhdl renameroo for output signals
  pcp_cpu_instruction_master_requests_cfi_flash_0_s1 <= internal_pcp_cpu_instruction_master_requests_cfi_flash_0_s1;
--synthesis translate_off
    --DBC3C40_SRAM_0/avalon_tristate_slave enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --incoming_tri_state_bridge_0_data_bit_0_is_x x check, which is an e_assign_is_x
    incoming_tri_state_bridge_0_data_bit_0_is_x <= A_WE_StdLogic(is_x(std_ulogic(internal_incoming_tri_state_bridge_0_data(0))), '1','0');
    --Crush incoming_tri_state_bridge_0_data_with_Xs_converted_to_0[0] Xs to 0, which is an e_assign
    incoming_tri_state_bridge_0_data_with_Xs_converted_to_0(0) <= A_WE_StdLogic((std_logic'(incoming_tri_state_bridge_0_data_bit_0_is_x) = '1'), std_logic'('0'), internal_incoming_tri_state_bridge_0_data(0));
    --incoming_tri_state_bridge_0_data_bit_1_is_x x check, which is an e_assign_is_x
    incoming_tri_state_bridge_0_data_bit_1_is_x <= A_WE_StdLogic(is_x(std_ulogic(internal_incoming_tri_state_bridge_0_data(1))), '1','0');
    --Crush incoming_tri_state_bridge_0_data_with_Xs_converted_to_0[1] Xs to 0, which is an e_assign
    incoming_tri_state_bridge_0_data_with_Xs_converted_to_0(1) <= A_WE_StdLogic((std_logic'(incoming_tri_state_bridge_0_data_bit_1_is_x) = '1'), std_logic'('0'), internal_incoming_tri_state_bridge_0_data(1));
    --incoming_tri_state_bridge_0_data_bit_2_is_x x check, which is an e_assign_is_x
    incoming_tri_state_bridge_0_data_bit_2_is_x <= A_WE_StdLogic(is_x(std_ulogic(internal_incoming_tri_state_bridge_0_data(2))), '1','0');
    --Crush incoming_tri_state_bridge_0_data_with_Xs_converted_to_0[2] Xs to 0, which is an e_assign
    incoming_tri_state_bridge_0_data_with_Xs_converted_to_0(2) <= A_WE_StdLogic((std_logic'(incoming_tri_state_bridge_0_data_bit_2_is_x) = '1'), std_logic'('0'), internal_incoming_tri_state_bridge_0_data(2));
    --incoming_tri_state_bridge_0_data_bit_3_is_x x check, which is an e_assign_is_x
    incoming_tri_state_bridge_0_data_bit_3_is_x <= A_WE_StdLogic(is_x(std_ulogic(internal_incoming_tri_state_bridge_0_data(3))), '1','0');
    --Crush incoming_tri_state_bridge_0_data_with_Xs_converted_to_0[3] Xs to 0, which is an e_assign
    incoming_tri_state_bridge_0_data_with_Xs_converted_to_0(3) <= A_WE_StdLogic((std_logic'(incoming_tri_state_bridge_0_data_bit_3_is_x) = '1'), std_logic'('0'), internal_incoming_tri_state_bridge_0_data(3));
    --incoming_tri_state_bridge_0_data_bit_4_is_x x check, which is an e_assign_is_x
    incoming_tri_state_bridge_0_data_bit_4_is_x <= A_WE_StdLogic(is_x(std_ulogic(internal_incoming_tri_state_bridge_0_data(4))), '1','0');
    --Crush incoming_tri_state_bridge_0_data_with_Xs_converted_to_0[4] Xs to 0, which is an e_assign
    incoming_tri_state_bridge_0_data_with_Xs_converted_to_0(4) <= A_WE_StdLogic((std_logic'(incoming_tri_state_bridge_0_data_bit_4_is_x) = '1'), std_logic'('0'), internal_incoming_tri_state_bridge_0_data(4));
    --incoming_tri_state_bridge_0_data_bit_5_is_x x check, which is an e_assign_is_x
    incoming_tri_state_bridge_0_data_bit_5_is_x <= A_WE_StdLogic(is_x(std_ulogic(internal_incoming_tri_state_bridge_0_data(5))), '1','0');
    --Crush incoming_tri_state_bridge_0_data_with_Xs_converted_to_0[5] Xs to 0, which is an e_assign
    incoming_tri_state_bridge_0_data_with_Xs_converted_to_0(5) <= A_WE_StdLogic((std_logic'(incoming_tri_state_bridge_0_data_bit_5_is_x) = '1'), std_logic'('0'), internal_incoming_tri_state_bridge_0_data(5));
    --incoming_tri_state_bridge_0_data_bit_6_is_x x check, which is an e_assign_is_x
    incoming_tri_state_bridge_0_data_bit_6_is_x <= A_WE_StdLogic(is_x(std_ulogic(internal_incoming_tri_state_bridge_0_data(6))), '1','0');
    --Crush incoming_tri_state_bridge_0_data_with_Xs_converted_to_0[6] Xs to 0, which is an e_assign
    incoming_tri_state_bridge_0_data_with_Xs_converted_to_0(6) <= A_WE_StdLogic((std_logic'(incoming_tri_state_bridge_0_data_bit_6_is_x) = '1'), std_logic'('0'), internal_incoming_tri_state_bridge_0_data(6));
    --incoming_tri_state_bridge_0_data_bit_7_is_x x check, which is an e_assign_is_x
    incoming_tri_state_bridge_0_data_bit_7_is_x <= A_WE_StdLogic(is_x(std_ulogic(internal_incoming_tri_state_bridge_0_data(7))), '1','0');
    --Crush incoming_tri_state_bridge_0_data_with_Xs_converted_to_0[7] Xs to 0, which is an e_assign
    incoming_tri_state_bridge_0_data_with_Xs_converted_to_0(7) <= A_WE_StdLogic((std_logic'(incoming_tri_state_bridge_0_data_bit_7_is_x) = '1'), std_logic'('0'), internal_incoming_tri_state_bridge_0_data(7));
    --incoming_tri_state_bridge_0_data_bit_8_is_x x check, which is an e_assign_is_x
    incoming_tri_state_bridge_0_data_bit_8_is_x <= A_WE_StdLogic(is_x(std_ulogic(internal_incoming_tri_state_bridge_0_data(8))), '1','0');
    --Crush incoming_tri_state_bridge_0_data_with_Xs_converted_to_0[8] Xs to 0, which is an e_assign
    incoming_tri_state_bridge_0_data_with_Xs_converted_to_0(8) <= A_WE_StdLogic((std_logic'(incoming_tri_state_bridge_0_data_bit_8_is_x) = '1'), std_logic'('0'), internal_incoming_tri_state_bridge_0_data(8));
    --incoming_tri_state_bridge_0_data_bit_9_is_x x check, which is an e_assign_is_x
    incoming_tri_state_bridge_0_data_bit_9_is_x <= A_WE_StdLogic(is_x(std_ulogic(internal_incoming_tri_state_bridge_0_data(9))), '1','0');
    --Crush incoming_tri_state_bridge_0_data_with_Xs_converted_to_0[9] Xs to 0, which is an e_assign
    incoming_tri_state_bridge_0_data_with_Xs_converted_to_0(9) <= A_WE_StdLogic((std_logic'(incoming_tri_state_bridge_0_data_bit_9_is_x) = '1'), std_logic'('0'), internal_incoming_tri_state_bridge_0_data(9));
    --incoming_tri_state_bridge_0_data_bit_10_is_x x check, which is an e_assign_is_x
    incoming_tri_state_bridge_0_data_bit_10_is_x <= A_WE_StdLogic(is_x(std_ulogic(internal_incoming_tri_state_bridge_0_data(10))), '1','0');
    --Crush incoming_tri_state_bridge_0_data_with_Xs_converted_to_0[10] Xs to 0, which is an e_assign
    incoming_tri_state_bridge_0_data_with_Xs_converted_to_0(10) <= A_WE_StdLogic((std_logic'(incoming_tri_state_bridge_0_data_bit_10_is_x) = '1'), std_logic'('0'), internal_incoming_tri_state_bridge_0_data(10));
    --incoming_tri_state_bridge_0_data_bit_11_is_x x check, which is an e_assign_is_x
    incoming_tri_state_bridge_0_data_bit_11_is_x <= A_WE_StdLogic(is_x(std_ulogic(internal_incoming_tri_state_bridge_0_data(11))), '1','0');
    --Crush incoming_tri_state_bridge_0_data_with_Xs_converted_to_0[11] Xs to 0, which is an e_assign
    incoming_tri_state_bridge_0_data_with_Xs_converted_to_0(11) <= A_WE_StdLogic((std_logic'(incoming_tri_state_bridge_0_data_bit_11_is_x) = '1'), std_logic'('0'), internal_incoming_tri_state_bridge_0_data(11));
    --incoming_tri_state_bridge_0_data_bit_12_is_x x check, which is an e_assign_is_x
    incoming_tri_state_bridge_0_data_bit_12_is_x <= A_WE_StdLogic(is_x(std_ulogic(internal_incoming_tri_state_bridge_0_data(12))), '1','0');
    --Crush incoming_tri_state_bridge_0_data_with_Xs_converted_to_0[12] Xs to 0, which is an e_assign
    incoming_tri_state_bridge_0_data_with_Xs_converted_to_0(12) <= A_WE_StdLogic((std_logic'(incoming_tri_state_bridge_0_data_bit_12_is_x) = '1'), std_logic'('0'), internal_incoming_tri_state_bridge_0_data(12));
    --incoming_tri_state_bridge_0_data_bit_13_is_x x check, which is an e_assign_is_x
    incoming_tri_state_bridge_0_data_bit_13_is_x <= A_WE_StdLogic(is_x(std_ulogic(internal_incoming_tri_state_bridge_0_data(13))), '1','0');
    --Crush incoming_tri_state_bridge_0_data_with_Xs_converted_to_0[13] Xs to 0, which is an e_assign
    incoming_tri_state_bridge_0_data_with_Xs_converted_to_0(13) <= A_WE_StdLogic((std_logic'(incoming_tri_state_bridge_0_data_bit_13_is_x) = '1'), std_logic'('0'), internal_incoming_tri_state_bridge_0_data(13));
    --incoming_tri_state_bridge_0_data_bit_14_is_x x check, which is an e_assign_is_x
    incoming_tri_state_bridge_0_data_bit_14_is_x <= A_WE_StdLogic(is_x(std_ulogic(internal_incoming_tri_state_bridge_0_data(14))), '1','0');
    --Crush incoming_tri_state_bridge_0_data_with_Xs_converted_to_0[14] Xs to 0, which is an e_assign
    incoming_tri_state_bridge_0_data_with_Xs_converted_to_0(14) <= A_WE_StdLogic((std_logic'(incoming_tri_state_bridge_0_data_bit_14_is_x) = '1'), std_logic'('0'), internal_incoming_tri_state_bridge_0_data(14));
    --incoming_tri_state_bridge_0_data_bit_15_is_x x check, which is an e_assign_is_x
    incoming_tri_state_bridge_0_data_bit_15_is_x <= A_WE_StdLogic(is_x(std_ulogic(internal_incoming_tri_state_bridge_0_data(15))), '1','0');
    --Crush incoming_tri_state_bridge_0_data_with_Xs_converted_to_0[15] Xs to 0, which is an e_assign
    incoming_tri_state_bridge_0_data_with_Xs_converted_to_0(15) <= A_WE_StdLogic((std_logic'(incoming_tri_state_bridge_0_data_bit_15_is_x) = '1'), std_logic'('0'), internal_incoming_tri_state_bridge_0_data(15));
    --cfi_flash_0/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --grant signals are active simultaneously, which is an e_process
    process (clk)
    VARIABLE write_line51 : line;
    begin
      if clk'event and clk = '1' then
        if (std_logic_vector'("0000000000000000000000000000") & (((std_logic_vector'("0") & (((std_logic_vector'("0") & (((std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(internal_pcp_cpu_data_master_granted_DBC3C40_SRAM_0_avalon_tristate_slave))) + (std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(internal_pcp_cpu_data_master_granted_cfi_flash_0_s1)))))) + (std_logic_vector'("00") & (A_TOSTDLOGICVECTOR(internal_pcp_cpu_instruction_master_granted_DBC3C40_SRAM_0_avalon_tristate_slave)))))) + (std_logic_vector'("000") & (A_TOSTDLOGICVECTOR(internal_pcp_cpu_instruction_master_granted_cfi_flash_0_s1))))))>std_logic_vector'("00000000000000000000000000000001") then 
          write(write_line51, now);
          write(write_line51, string'(": "));
          write(write_line51, string'("> 1 of grant signals are active simultaneously"));
          write(output, write_line51.all);
          deallocate (write_line51);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --saved_grant signals are active simultaneously, which is an e_process
    process (clk)
    VARIABLE write_line52 : line;
    begin
      if clk'event and clk = '1' then
        if (std_logic_vector'("0000000000000000000000000000") & (((std_logic_vector'("0") & (((std_logic_vector'("0") & (((std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(pcp_cpu_data_master_saved_grant_DBC3C40_SRAM_0_avalon_tristate_slave))) + (std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(pcp_cpu_data_master_saved_grant_cfi_flash_0_s1)))))) + (std_logic_vector'("00") & (A_TOSTDLOGICVECTOR(pcp_cpu_instruction_master_saved_grant_DBC3C40_SRAM_0_avalon_tristate_slave)))))) + (std_logic_vector'("000") & (A_TOSTDLOGICVECTOR(pcp_cpu_instruction_master_saved_grant_cfi_flash_0_s1))))))>std_logic_vector'("00000000000000000000000000000001") then 
          write(write_line52, now);
          write(write_line52, string'(": "));
          write(write_line52, string'("> 1 of saved_grant signals are active simultaneously"));
          write(output, write_line52.all);
          deallocate (write_line52);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on
--synthesis read_comments_as_HDL on
--    
--    incoming_tri_state_bridge_0_data_with_Xs_converted_to_0 <= internal_incoming_tri_state_bridge_0_data;
--synthesis read_comments_as_HDL off

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity tri_state_bridge_0_bridge_arbitrator is 
end entity tri_state_bridge_0_bridge_arbitrator;


architecture europa of tri_state_bridge_0_bridge_arbitrator is

begin


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity niosII_openMac_reset_clk50Meg_domain_synch_module is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC
              );
end entity niosII_openMac_reset_clk50Meg_domain_synch_module;


architecture europa of niosII_openMac_reset_clk50Meg_domain_synch_module is
                signal data_in_d1 :  STD_LOGIC;
attribute ALTERA_ATTRIBUTE : string;
attribute ALTERA_ATTRIBUTE of data_in_d1 : signal is "{-from ""*""} CUT=ON ; PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101";
attribute ALTERA_ATTRIBUTE of data_out : signal is "PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101";

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      data_in_d1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      data_in_d1 <= data_in;
    end if;

  end process;

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      data_out <= std_logic'('0');
    elsif clk'event and clk = '1' then
      data_out <= data_in_d1;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity niosII_openMac_reset_clk90Meg_domain_synch_module is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC
              );
end entity niosII_openMac_reset_clk90Meg_domain_synch_module;


architecture europa of niosII_openMac_reset_clk90Meg_domain_synch_module is
                signal data_in_d1 :  STD_LOGIC;
attribute ALTERA_ATTRIBUTE : string;
attribute ALTERA_ATTRIBUTE of data_in_d1 : signal is "{-from ""*""} CUT=ON ; PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101";
attribute ALTERA_ATTRIBUTE of data_out : signal is "PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101";

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      data_in_d1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      data_in_d1 <= data_in;
    end if;

  end process;

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      data_out <= std_logic'('0');
    elsif clk'event and clk = '1' then
      data_out <= data_in_d1;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity niosII_openMac_reset_clk_0_domain_synch_module is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC
              );
end entity niosII_openMac_reset_clk_0_domain_synch_module;


architecture europa of niosII_openMac_reset_clk_0_domain_synch_module is
                signal data_in_d1 :  STD_LOGIC;
attribute ALTERA_ATTRIBUTE : string;
attribute ALTERA_ATTRIBUTE of data_in_d1 : signal is "{-from ""*""} CUT=ON ; PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101";
attribute ALTERA_ATTRIBUTE of data_out : signal is "PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101";

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      data_in_d1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      data_in_d1 <= data_in;
    end if;

  end process;

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      data_out <= std_logic'('0');
    elsif clk'event and clk = '1' then
      data_out <= data_in_d1;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity niosII_openMac_reset_clk25Meg_domain_synch_module is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC
              );
end entity niosII_openMac_reset_clk25Meg_domain_synch_module;


architecture europa of niosII_openMac_reset_clk25Meg_domain_synch_module is
                signal data_in_d1 :  STD_LOGIC;
attribute ALTERA_ATTRIBUTE : string;
attribute ALTERA_ATTRIBUTE of data_in_d1 : signal is "{-from ""*""} CUT=ON ; PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101";
attribute ALTERA_ATTRIBUTE of data_out : signal is "PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101";

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      data_in_d1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      data_in_d1 <= data_in;
    end if;

  end process;

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      data_out <= std_logic'('0');
    elsif clk'event and clk = '1' then
      data_out <= data_in_d1;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity niosII_openMac is 
        port (
              -- 1) global signals:
                 signal clk100Meg180 : OUT STD_LOGIC;
                 signal clk25Meg : OUT STD_LOGIC;
                 signal clk50Meg : OUT STD_LOGIC;
                 signal clk90Meg : OUT STD_LOGIC;
                 signal clk90MegSDRAM : OUT STD_LOGIC;
                 signal clk_0 : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- the_OpenMAC_0
                 signal mii_Clk_from_the_OpenMAC_0 : OUT STD_LOGIC;
                 signal mii_Di_to_the_OpenMAC_0 : IN STD_LOGIC;
                 signal mii_Do_from_the_OpenMAC_0 : OUT STD_LOGIC;
                 signal mii_Doe_from_the_OpenMAC_0 : OUT STD_LOGIC;
                 signal mii_nResetOut_from_the_OpenMAC_0 : OUT STD_LOGIC;
                 signal rCrs_Dv_0_to_the_OpenMAC_0 : IN STD_LOGIC;
                 signal rCrs_Dv_1_to_the_OpenMAC_0 : IN STD_LOGIC;
                 signal rRx_Dat_0_to_the_OpenMAC_0 : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal rRx_Dat_1_to_the_OpenMAC_0 : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal rTx_Dat_0_from_the_OpenMAC_0 : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal rTx_Dat_1_from_the_OpenMAC_0 : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal rTx_En_0_from_the_OpenMAC_0 : OUT STD_LOGIC;
                 signal rTx_En_1_from_the_OpenMAC_0 : OUT STD_LOGIC;

              -- the_altpll_0
                 signal locked_from_the_altpll_0 : OUT STD_LOGIC;
                 signal phasedone_from_the_altpll_0 : OUT STD_LOGIC;

              -- the_button_pio
                 signal in_port_to_the_button_pio : IN STD_LOGIC_VECTOR (7 DOWNTO 0);

              -- the_digio_pio
                 signal bidir_port_to_and_from_the_digio_pio : INOUT STD_LOGIC_VECTOR (31 DOWNTO 0);

              -- the_epcs_flash_controller_0
                 signal data0_to_the_epcs_flash_controller_0 : IN STD_LOGIC;
                 signal dclk_from_the_epcs_flash_controller_0 : OUT STD_LOGIC;
                 signal sce_from_the_epcs_flash_controller_0 : OUT STD_LOGIC;
                 signal sdo_from_the_epcs_flash_controller_0 : OUT STD_LOGIC;

              -- the_irq_gen
                 signal out_port_from_the_irq_gen : OUT STD_LOGIC;

              -- the_node_switch_pio
                 signal in_port_to_the_node_switch_pio : IN STD_LOGIC_VECTOR (7 DOWNTO 0);

              -- the_portconf_pio
                 signal in_port_to_the_portconf_pio : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal out_port_from_the_portconf_pio : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);

              -- the_sdram_0
                 signal zs_addr_from_the_sdram_0 : OUT STD_LOGIC_VECTOR (11 DOWNTO 0);
                 signal zs_ba_from_the_sdram_0 : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal zs_cas_n_from_the_sdram_0 : OUT STD_LOGIC;
                 signal zs_cke_from_the_sdram_0 : OUT STD_LOGIC;
                 signal zs_cs_n_from_the_sdram_0 : OUT STD_LOGIC;
                 signal zs_dq_to_and_from_the_sdram_0 : INOUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal zs_dqm_from_the_sdram_0 : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal zs_ras_n_from_the_sdram_0 : OUT STD_LOGIC;
                 signal zs_we_n_from_the_sdram_0 : OUT STD_LOGIC;

              -- the_status_led_pio
                 signal out_port_from_the_status_led_pio : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);

              -- the_sync_irq
                 signal in_port_to_the_sync_irq : IN STD_LOGIC;

              -- the_tri_state_bridge_0_avalon_slave
                 signal ben_to_the_DBC3C40_SRAM_0 : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal ncs_to_the_DBC3C40_SRAM_0 : OUT STD_LOGIC;
                 signal select_n_to_the_cfi_flash_0 : OUT STD_LOGIC;
                 signal tri_state_bridge_0_address : OUT STD_LOGIC_VECTOR (22 DOWNTO 0);
                 signal tri_state_bridge_0_data : INOUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal tri_state_bridge_0_readn : OUT STD_LOGIC;
                 signal tri_state_bridge_0_writen : OUT STD_LOGIC
              );
end entity niosII_openMac;


architecture europa of niosII_openMac is
component OpenMAC_0_CMP_arbitrator is 
           port (
                 -- inputs:
                    signal OpenMAC_0_CMP_irq : IN STD_LOGIC;
                    signal OpenMAC_0_CMP_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal clk : IN STD_LOGIC;
                    signal niosII_openMac_clock_1_out_address_to_slave : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal niosII_openMac_clock_1_out_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal niosII_openMac_clock_1_out_read : IN STD_LOGIC;
                    signal niosII_openMac_clock_1_out_write : IN STD_LOGIC;
                    signal niosII_openMac_clock_1_out_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal OpenMAC_0_CMP_address : OUT STD_LOGIC;
                    signal OpenMAC_0_CMP_byteenable_n : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal OpenMAC_0_CMP_chipselect : OUT STD_LOGIC;
                    signal OpenMAC_0_CMP_irq_from_sa : OUT STD_LOGIC;
                    signal OpenMAC_0_CMP_read_n : OUT STD_LOGIC;
                    signal OpenMAC_0_CMP_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal OpenMAC_0_CMP_reset_n : OUT STD_LOGIC;
                    signal OpenMAC_0_CMP_write_n : OUT STD_LOGIC;
                    signal OpenMAC_0_CMP_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal d1_OpenMAC_0_CMP_end_xfer : OUT STD_LOGIC;
                    signal niosII_openMac_clock_1_out_granted_OpenMAC_0_CMP : OUT STD_LOGIC;
                    signal niosII_openMac_clock_1_out_qualified_request_OpenMAC_0_CMP : OUT STD_LOGIC;
                    signal niosII_openMac_clock_1_out_read_data_valid_OpenMAC_0_CMP : OUT STD_LOGIC;
                    signal niosII_openMac_clock_1_out_requests_OpenMAC_0_CMP : OUT STD_LOGIC
                 );
end component OpenMAC_0_CMP_arbitrator;

component OpenMAC_0_REG_arbitrator is 
           port (
                 -- inputs:
                    signal OpenMAC_0_REG_irq : IN STD_LOGIC;
                    signal OpenMAC_0_REG_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal clk : IN STD_LOGIC;
                    signal niosII_openMac_clock_2_out_address_to_slave : IN STD_LOGIC_VECTOR (12 DOWNTO 0);
                    signal niosII_openMac_clock_2_out_byteenable : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal niosII_openMac_clock_2_out_read : IN STD_LOGIC;
                    signal niosII_openMac_clock_2_out_write : IN STD_LOGIC;
                    signal niosII_openMac_clock_2_out_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal OpenMAC_0_REG_address : OUT STD_LOGIC_VECTOR (11 DOWNTO 0);
                    signal OpenMAC_0_REG_byteenable_n : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal OpenMAC_0_REG_chipselect : OUT STD_LOGIC;
                    signal OpenMAC_0_REG_irq_from_sa : OUT STD_LOGIC;
                    signal OpenMAC_0_REG_read_n : OUT STD_LOGIC;
                    signal OpenMAC_0_REG_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal OpenMAC_0_REG_write_n : OUT STD_LOGIC;
                    signal OpenMAC_0_REG_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal d1_OpenMAC_0_REG_end_xfer : OUT STD_LOGIC;
                    signal niosII_openMac_clock_2_out_granted_OpenMAC_0_REG : OUT STD_LOGIC;
                    signal niosII_openMac_clock_2_out_qualified_request_OpenMAC_0_REG : OUT STD_LOGIC;
                    signal niosII_openMac_clock_2_out_read_data_valid_OpenMAC_0_REG : OUT STD_LOGIC;
                    signal niosII_openMac_clock_2_out_requests_OpenMAC_0_REG : OUT STD_LOGIC
                 );
end component OpenMAC_0_REG_arbitrator;

component OpenMAC_0_iBuf_arbitrator is 
           port (
                 -- inputs:
                    signal OpenMAC_0_iBuf_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal clk : IN STD_LOGIC;
                    signal pcp_cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (25 DOWNTO 0);
                    signal pcp_cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal pcp_cpu_data_master_read : IN STD_LOGIC;
                    signal pcp_cpu_data_master_waitrequest : IN STD_LOGIC;
                    signal pcp_cpu_data_master_write : IN STD_LOGIC;
                    signal pcp_cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal OpenMAC_0_iBuf_address : OUT STD_LOGIC_VECTOR (12 DOWNTO 0);
                    signal OpenMAC_0_iBuf_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal OpenMAC_0_iBuf_chipselect : OUT STD_LOGIC;
                    signal OpenMAC_0_iBuf_read_n : OUT STD_LOGIC;
                    signal OpenMAC_0_iBuf_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal OpenMAC_0_iBuf_wait_counter_eq_0 : OUT STD_LOGIC;
                    signal OpenMAC_0_iBuf_write_n : OUT STD_LOGIC;
                    signal OpenMAC_0_iBuf_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal d1_OpenMAC_0_iBuf_end_xfer : OUT STD_LOGIC;
                    signal pcp_cpu_data_master_granted_OpenMAC_0_iBuf : OUT STD_LOGIC;
                    signal pcp_cpu_data_master_qualified_request_OpenMAC_0_iBuf : OUT STD_LOGIC;
                    signal pcp_cpu_data_master_read_data_valid_OpenMAC_0_iBuf : OUT STD_LOGIC;
                    signal pcp_cpu_data_master_requests_OpenMAC_0_iBuf : OUT STD_LOGIC
                 );
end component OpenMAC_0_iBuf_arbitrator;

component OpenMAC_0 is 
           port (
                 -- inputs:
                    signal Clk50 : IN STD_LOGIC;
                    signal ClkFaster : IN STD_LOGIC;
                    signal Reset_n : IN STD_LOGIC;
                    signal iBuf_address : IN STD_LOGIC_VECTOR (12 DOWNTO 0);
                    signal iBuf_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal iBuf_chipselect : IN STD_LOGIC;
                    signal iBuf_read_n : IN STD_LOGIC;
                    signal iBuf_write_n : IN STD_LOGIC;
                    signal iBuf_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal mii_Di : IN STD_LOGIC;
                    signal rCrs_Dv_0 : IN STD_LOGIC;
                    signal rCrs_Dv_1 : IN STD_LOGIC;
                    signal rRx_Dat_0 : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal rRx_Dat_1 : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal s_address : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
                    signal s_byteenable_n : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal s_chipselect : IN STD_LOGIC;
                    signal s_read_n : IN STD_LOGIC;
                    signal s_write_n : IN STD_LOGIC;
                    signal s_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal t_address : IN STD_LOGIC_VECTOR (0 DOWNTO 0);
                    signal t_byteenable_n : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal t_chipselect : IN STD_LOGIC;
                    signal t_read_n : IN STD_LOGIC;
                    signal t_write_n : IN STD_LOGIC;
                    signal t_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal iBuf_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal mii_Clk : OUT STD_LOGIC;
                    signal mii_Do : OUT STD_LOGIC;
                    signal mii_Doe : OUT STD_LOGIC;
                    signal mii_nResetOut : OUT STD_LOGIC;
                    signal rTx_Dat_0 : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal rTx_Dat_1 : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal rTx_En_0 : OUT STD_LOGIC;
                    signal rTx_En_1 : OUT STD_LOGIC;
                    signal s_IRQ : OUT STD_LOGIC;
                    signal s_readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal t_IRQ : OUT STD_LOGIC;
                    signal t_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
                 );
end component OpenMAC_0;

component altpll_0_pll_slave_arbitrator is 
           port (
                 -- inputs:
                    signal altpll_0_pll_slave_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal clk : IN STD_LOGIC;
                    signal niosII_openMac_clock_3_out_address_to_slave : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal niosII_openMac_clock_3_out_read : IN STD_LOGIC;
                    signal niosII_openMac_clock_3_out_write : IN STD_LOGIC;
                    signal niosII_openMac_clock_3_out_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal altpll_0_pll_slave_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal altpll_0_pll_slave_read : OUT STD_LOGIC;
                    signal altpll_0_pll_slave_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal altpll_0_pll_slave_reset : OUT STD_LOGIC;
                    signal altpll_0_pll_slave_write : OUT STD_LOGIC;
                    signal altpll_0_pll_slave_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal d1_altpll_0_pll_slave_end_xfer : OUT STD_LOGIC;
                    signal niosII_openMac_clock_3_out_granted_altpll_0_pll_slave : OUT STD_LOGIC;
                    signal niosII_openMac_clock_3_out_qualified_request_altpll_0_pll_slave : OUT STD_LOGIC;
                    signal niosII_openMac_clock_3_out_read_data_valid_altpll_0_pll_slave : OUT STD_LOGIC;
                    signal niosII_openMac_clock_3_out_requests_altpll_0_pll_slave : OUT STD_LOGIC
                 );
end component altpll_0_pll_slave_arbitrator;

component altpll_0 is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal clk : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal c0 : OUT STD_LOGIC;
                    signal c1 : OUT STD_LOGIC;
                    signal c2 : OUT STD_LOGIC;
                    signal c3 : OUT STD_LOGIC;
                    signal c4 : OUT STD_LOGIC;
                    signal locked : OUT STD_LOGIC;
                    signal phasedone : OUT STD_LOGIC;
                    signal readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
                 );
end component altpll_0;

component ap_cpu_jtag_debug_module_arbitrator is 
           port (
                 -- inputs:
                    signal ap_cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (25 DOWNTO 0);
                    signal ap_cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal ap_cpu_data_master_debugaccess : IN STD_LOGIC;
                    signal ap_cpu_data_master_read : IN STD_LOGIC;
                    signal ap_cpu_data_master_waitrequest : IN STD_LOGIC;
                    signal ap_cpu_data_master_write : IN STD_LOGIC;
                    signal ap_cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal ap_cpu_instruction_master_address_to_slave : IN STD_LOGIC_VECTOR (25 DOWNTO 0);
                    signal ap_cpu_instruction_master_latency_counter : IN STD_LOGIC;
                    signal ap_cpu_instruction_master_read : IN STD_LOGIC;
                    signal ap_cpu_instruction_master_read_data_valid_sdram_0_s1_shift_register : IN STD_LOGIC;
                    signal ap_cpu_jtag_debug_module_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal ap_cpu_jtag_debug_module_resetrequest : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal ap_cpu_data_master_granted_ap_cpu_jtag_debug_module : OUT STD_LOGIC;
                    signal ap_cpu_data_master_qualified_request_ap_cpu_jtag_debug_module : OUT STD_LOGIC;
                    signal ap_cpu_data_master_read_data_valid_ap_cpu_jtag_debug_module : OUT STD_LOGIC;
                    signal ap_cpu_data_master_requests_ap_cpu_jtag_debug_module : OUT STD_LOGIC;
                    signal ap_cpu_instruction_master_granted_ap_cpu_jtag_debug_module : OUT STD_LOGIC;
                    signal ap_cpu_instruction_master_qualified_request_ap_cpu_jtag_debug_module : OUT STD_LOGIC;
                    signal ap_cpu_instruction_master_read_data_valid_ap_cpu_jtag_debug_module : OUT STD_LOGIC;
                    signal ap_cpu_instruction_master_requests_ap_cpu_jtag_debug_module : OUT STD_LOGIC;
                    signal ap_cpu_jtag_debug_module_address : OUT STD_LOGIC_VECTOR (8 DOWNTO 0);
                    signal ap_cpu_jtag_debug_module_begintransfer : OUT STD_LOGIC;
                    signal ap_cpu_jtag_debug_module_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal ap_cpu_jtag_debug_module_chipselect : OUT STD_LOGIC;
                    signal ap_cpu_jtag_debug_module_debugaccess : OUT STD_LOGIC;
                    signal ap_cpu_jtag_debug_module_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal ap_cpu_jtag_debug_module_reset_n : OUT STD_LOGIC;
                    signal ap_cpu_jtag_debug_module_resetrequest_from_sa : OUT STD_LOGIC;
                    signal ap_cpu_jtag_debug_module_write : OUT STD_LOGIC;
                    signal ap_cpu_jtag_debug_module_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal d1_ap_cpu_jtag_debug_module_end_xfer : OUT STD_LOGIC
                 );
end component ap_cpu_jtag_debug_module_arbitrator;

component ap_cpu_data_master_arbitrator is 
           port (
                 -- inputs:
                    signal ap_cpu_data_master_address : IN STD_LOGIC_VECTOR (25 DOWNTO 0);
                    signal ap_cpu_data_master_granted_ap_cpu_jtag_debug_module : IN STD_LOGIC;
                    signal ap_cpu_data_master_granted_clock_crossing_1_s1 : IN STD_LOGIC;
                    signal ap_cpu_data_master_granted_cnApi_Av2Av_0_ap : IN STD_LOGIC;
                    signal ap_cpu_data_master_granted_jtag_uart_1_avalon_jtag_slave : IN STD_LOGIC;
                    signal ap_cpu_data_master_granted_sdram_0_s1 : IN STD_LOGIC;
                    signal ap_cpu_data_master_qualified_request_ap_cpu_jtag_debug_module : IN STD_LOGIC;
                    signal ap_cpu_data_master_qualified_request_clock_crossing_1_s1 : IN STD_LOGIC;
                    signal ap_cpu_data_master_qualified_request_cnApi_Av2Av_0_ap : IN STD_LOGIC;
                    signal ap_cpu_data_master_qualified_request_jtag_uart_1_avalon_jtag_slave : IN STD_LOGIC;
                    signal ap_cpu_data_master_qualified_request_sdram_0_s1 : IN STD_LOGIC;
                    signal ap_cpu_data_master_read : IN STD_LOGIC;
                    signal ap_cpu_data_master_read_data_valid_ap_cpu_jtag_debug_module : IN STD_LOGIC;
                    signal ap_cpu_data_master_read_data_valid_clock_crossing_1_s1 : IN STD_LOGIC;
                    signal ap_cpu_data_master_read_data_valid_clock_crossing_1_s1_shift_register : IN STD_LOGIC;
                    signal ap_cpu_data_master_read_data_valid_cnApi_Av2Av_0_ap : IN STD_LOGIC;
                    signal ap_cpu_data_master_read_data_valid_jtag_uart_1_avalon_jtag_slave : IN STD_LOGIC;
                    signal ap_cpu_data_master_read_data_valid_sdram_0_s1 : IN STD_LOGIC;
                    signal ap_cpu_data_master_read_data_valid_sdram_0_s1_shift_register : IN STD_LOGIC;
                    signal ap_cpu_data_master_requests_ap_cpu_jtag_debug_module : IN STD_LOGIC;
                    signal ap_cpu_data_master_requests_clock_crossing_1_s1 : IN STD_LOGIC;
                    signal ap_cpu_data_master_requests_cnApi_Av2Av_0_ap : IN STD_LOGIC;
                    signal ap_cpu_data_master_requests_jtag_uart_1_avalon_jtag_slave : IN STD_LOGIC;
                    signal ap_cpu_data_master_requests_sdram_0_s1 : IN STD_LOGIC;
                    signal ap_cpu_data_master_write : IN STD_LOGIC;
                    signal ap_cpu_jtag_debug_module_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal clk : IN STD_LOGIC;
                    signal clk90Meg : IN STD_LOGIC;
                    signal clk90Meg_reset_n : IN STD_LOGIC;
                    signal clock_crossing_1_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal clock_crossing_1_s1_waitrequest_from_sa : IN STD_LOGIC;
                    signal cnApi_Av2Av_0_ap_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal cnApi_Av2Av_0_ap_wait_counter_eq_0 : IN STD_LOGIC;
                    signal d1_ap_cpu_jtag_debug_module_end_xfer : IN STD_LOGIC;
                    signal d1_clock_crossing_1_s1_end_xfer : IN STD_LOGIC;
                    signal d1_cnApi_Av2Av_0_ap_end_xfer : IN STD_LOGIC;
                    signal d1_jtag_uart_1_avalon_jtag_slave_end_xfer : IN STD_LOGIC;
                    signal d1_sdram_0_s1_end_xfer : IN STD_LOGIC;
                    signal jtag_uart_1_avalon_jtag_slave_irq_from_sa : IN STD_LOGIC;
                    signal jtag_uart_1_avalon_jtag_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal jtag_uart_1_avalon_jtag_slave_waitrequest_from_sa : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sdram_0_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal sdram_0_s1_waitrequest_from_sa : IN STD_LOGIC;
                    signal sync_irq_s1_irq_from_sa : IN STD_LOGIC;
                    signal system_timer_ap_s1_irq_from_sa : IN STD_LOGIC;

                 -- outputs:
                    signal ap_cpu_data_master_address_to_slave : OUT STD_LOGIC_VECTOR (25 DOWNTO 0);
                    signal ap_cpu_data_master_irq : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal ap_cpu_data_master_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal ap_cpu_data_master_waitrequest : OUT STD_LOGIC
                 );
end component ap_cpu_data_master_arbitrator;

component ap_cpu_instruction_master_arbitrator is 
           port (
                 -- inputs:
                    signal ap_cpu_instruction_master_address : IN STD_LOGIC_VECTOR (25 DOWNTO 0);
                    signal ap_cpu_instruction_master_granted_ap_cpu_jtag_debug_module : IN STD_LOGIC;
                    signal ap_cpu_instruction_master_granted_sdram_0_s1 : IN STD_LOGIC;
                    signal ap_cpu_instruction_master_qualified_request_ap_cpu_jtag_debug_module : IN STD_LOGIC;
                    signal ap_cpu_instruction_master_qualified_request_sdram_0_s1 : IN STD_LOGIC;
                    signal ap_cpu_instruction_master_read : IN STD_LOGIC;
                    signal ap_cpu_instruction_master_read_data_valid_ap_cpu_jtag_debug_module : IN STD_LOGIC;
                    signal ap_cpu_instruction_master_read_data_valid_sdram_0_s1 : IN STD_LOGIC;
                    signal ap_cpu_instruction_master_read_data_valid_sdram_0_s1_shift_register : IN STD_LOGIC;
                    signal ap_cpu_instruction_master_requests_ap_cpu_jtag_debug_module : IN STD_LOGIC;
                    signal ap_cpu_instruction_master_requests_sdram_0_s1 : IN STD_LOGIC;
                    signal ap_cpu_jtag_debug_module_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal clk : IN STD_LOGIC;
                    signal d1_ap_cpu_jtag_debug_module_end_xfer : IN STD_LOGIC;
                    signal d1_sdram_0_s1_end_xfer : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sdram_0_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal sdram_0_s1_waitrequest_from_sa : IN STD_LOGIC;

                 -- outputs:
                    signal ap_cpu_instruction_master_address_to_slave : OUT STD_LOGIC_VECTOR (25 DOWNTO 0);
                    signal ap_cpu_instruction_master_latency_counter : OUT STD_LOGIC;
                    signal ap_cpu_instruction_master_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal ap_cpu_instruction_master_readdatavalid : OUT STD_LOGIC;
                    signal ap_cpu_instruction_master_waitrequest : OUT STD_LOGIC
                 );
end component ap_cpu_instruction_master_arbitrator;

component ap_cpu is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal d_irq : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal d_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal d_waitrequest : IN STD_LOGIC;
                    signal i_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal i_readdatavalid : IN STD_LOGIC;
                    signal i_waitrequest : IN STD_LOGIC;
                    signal jtag_debug_module_address : IN STD_LOGIC_VECTOR (8 DOWNTO 0);
                    signal jtag_debug_module_begintransfer : IN STD_LOGIC;
                    signal jtag_debug_module_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal jtag_debug_module_debugaccess : IN STD_LOGIC;
                    signal jtag_debug_module_select : IN STD_LOGIC;
                    signal jtag_debug_module_write : IN STD_LOGIC;
                    signal jtag_debug_module_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal d_address : OUT STD_LOGIC_VECTOR (25 DOWNTO 0);
                    signal d_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal d_read : OUT STD_LOGIC;
                    signal d_write : OUT STD_LOGIC;
                    signal d_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal i_address : OUT STD_LOGIC_VECTOR (25 DOWNTO 0);
                    signal i_read : OUT STD_LOGIC;
                    signal jtag_debug_module_debugaccess_to_roms : OUT STD_LOGIC;
                    signal jtag_debug_module_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal jtag_debug_module_resetrequest : OUT STD_LOGIC
                 );
end component ap_cpu;

component button_pio_s1_arbitrator is 
           port (
                 -- inputs:
                    signal button_pio_s1_readdata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal clk : IN STD_LOGIC;
                    signal clock_crossing_0_m1_address_to_slave : IN STD_LOGIC_VECTOR (6 DOWNTO 0);
                    signal clock_crossing_0_m1_latency_counter : IN STD_LOGIC;
                    signal clock_crossing_0_m1_nativeaddress : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
                    signal clock_crossing_0_m1_read : IN STD_LOGIC;
                    signal clock_crossing_0_m1_write : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal button_pio_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal button_pio_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal button_pio_s1_reset_n : OUT STD_LOGIC;
                    signal clock_crossing_0_m1_granted_button_pio_s1 : OUT STD_LOGIC;
                    signal clock_crossing_0_m1_qualified_request_button_pio_s1 : OUT STD_LOGIC;
                    signal clock_crossing_0_m1_read_data_valid_button_pio_s1 : OUT STD_LOGIC;
                    signal clock_crossing_0_m1_requests_button_pio_s1 : OUT STD_LOGIC;
                    signal d1_button_pio_s1_end_xfer : OUT STD_LOGIC
                 );
end component button_pio_s1_arbitrator;

component button_pio is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal clk : IN STD_LOGIC;
                    signal in_port : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal readdata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
                 );
end component button_pio;

component clock_crossing_0_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal clock_crossing_0_s1_endofpacket : IN STD_LOGIC;
                    signal clock_crossing_0_s1_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal clock_crossing_0_s1_readdatavalid : IN STD_LOGIC;
                    signal clock_crossing_0_s1_waitrequest : IN STD_LOGIC;
                    signal pcp_cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (25 DOWNTO 0);
                    signal pcp_cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal pcp_cpu_data_master_read : IN STD_LOGIC;
                    signal pcp_cpu_data_master_waitrequest : IN STD_LOGIC;
                    signal pcp_cpu_data_master_write : IN STD_LOGIC;
                    signal pcp_cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal clock_crossing_0_s1_address : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
                    signal clock_crossing_0_s1_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal clock_crossing_0_s1_endofpacket_from_sa : OUT STD_LOGIC;
                    signal clock_crossing_0_s1_nativeaddress : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
                    signal clock_crossing_0_s1_read : OUT STD_LOGIC;
                    signal clock_crossing_0_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal clock_crossing_0_s1_reset_n : OUT STD_LOGIC;
                    signal clock_crossing_0_s1_waitrequest_from_sa : OUT STD_LOGIC;
                    signal clock_crossing_0_s1_write : OUT STD_LOGIC;
                    signal clock_crossing_0_s1_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal d1_clock_crossing_0_s1_end_xfer : OUT STD_LOGIC;
                    signal pcp_cpu_data_master_granted_clock_crossing_0_s1 : OUT STD_LOGIC;
                    signal pcp_cpu_data_master_qualified_request_clock_crossing_0_s1 : OUT STD_LOGIC;
                    signal pcp_cpu_data_master_read_data_valid_clock_crossing_0_s1 : OUT STD_LOGIC;
                    signal pcp_cpu_data_master_read_data_valid_clock_crossing_0_s1_shift_register : OUT STD_LOGIC;
                    signal pcp_cpu_data_master_requests_clock_crossing_0_s1 : OUT STD_LOGIC
                 );
end component clock_crossing_0_s1_arbitrator;

component clock_crossing_0_m1_arbitrator is 
           port (
                 -- inputs:
                    signal button_pio_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal clk : IN STD_LOGIC;
                    signal clock_crossing_0_m1_address : IN STD_LOGIC_VECTOR (6 DOWNTO 0);
                    signal clock_crossing_0_m1_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal clock_crossing_0_m1_granted_button_pio_s1 : IN STD_LOGIC;
                    signal clock_crossing_0_m1_granted_irq_gen_s1 : IN STD_LOGIC;
                    signal clock_crossing_0_m1_granted_status_led_pio_s1 : IN STD_LOGIC;
                    signal clock_crossing_0_m1_granted_sysid_control_slave : IN STD_LOGIC;
                    signal clock_crossing_0_m1_granted_system_timer_s1 : IN STD_LOGIC;
                    signal clock_crossing_0_m1_qualified_request_button_pio_s1 : IN STD_LOGIC;
                    signal clock_crossing_0_m1_qualified_request_irq_gen_s1 : IN STD_LOGIC;
                    signal clock_crossing_0_m1_qualified_request_status_led_pio_s1 : IN STD_LOGIC;
                    signal clock_crossing_0_m1_qualified_request_sysid_control_slave : IN STD_LOGIC;
                    signal clock_crossing_0_m1_qualified_request_system_timer_s1 : IN STD_LOGIC;
                    signal clock_crossing_0_m1_read : IN STD_LOGIC;
                    signal clock_crossing_0_m1_read_data_valid_button_pio_s1 : IN STD_LOGIC;
                    signal clock_crossing_0_m1_read_data_valid_irq_gen_s1 : IN STD_LOGIC;
                    signal clock_crossing_0_m1_read_data_valid_status_led_pio_s1 : IN STD_LOGIC;
                    signal clock_crossing_0_m1_read_data_valid_sysid_control_slave : IN STD_LOGIC;
                    signal clock_crossing_0_m1_read_data_valid_system_timer_s1 : IN STD_LOGIC;
                    signal clock_crossing_0_m1_requests_button_pio_s1 : IN STD_LOGIC;
                    signal clock_crossing_0_m1_requests_irq_gen_s1 : IN STD_LOGIC;
                    signal clock_crossing_0_m1_requests_status_led_pio_s1 : IN STD_LOGIC;
                    signal clock_crossing_0_m1_requests_sysid_control_slave : IN STD_LOGIC;
                    signal clock_crossing_0_m1_requests_system_timer_s1 : IN STD_LOGIC;
                    signal clock_crossing_0_m1_write : IN STD_LOGIC;
                    signal clock_crossing_0_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal d1_button_pio_s1_end_xfer : IN STD_LOGIC;
                    signal d1_irq_gen_s1_end_xfer : IN STD_LOGIC;
                    signal d1_status_led_pio_s1_end_xfer : IN STD_LOGIC;
                    signal d1_sysid_control_slave_end_xfer : IN STD_LOGIC;
                    signal d1_system_timer_s1_end_xfer : IN STD_LOGIC;
                    signal irq_gen_s1_readdata_from_sa : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal status_led_pio_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal sysid_control_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal system_timer_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

                 -- outputs:
                    signal clock_crossing_0_m1_address_to_slave : OUT STD_LOGIC_VECTOR (6 DOWNTO 0);
                    signal clock_crossing_0_m1_latency_counter : OUT STD_LOGIC;
                    signal clock_crossing_0_m1_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal clock_crossing_0_m1_readdatavalid : OUT STD_LOGIC;
                    signal clock_crossing_0_m1_reset_n : OUT STD_LOGIC;
                    signal clock_crossing_0_m1_waitrequest : OUT STD_LOGIC
                 );
end component clock_crossing_0_m1_arbitrator;

component clock_crossing_0 is 
           port (
                 -- inputs:
                    signal master_clk : IN STD_LOGIC;
                    signal master_endofpacket : IN STD_LOGIC;
                    signal master_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal master_readdatavalid : IN STD_LOGIC;
                    signal master_reset_n : IN STD_LOGIC;
                    signal master_waitrequest : IN STD_LOGIC;
                    signal slave_address : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
                    signal slave_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal slave_clk : IN STD_LOGIC;
                    signal slave_nativeaddress : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
                    signal slave_read : IN STD_LOGIC;
                    signal slave_reset_n : IN STD_LOGIC;
                    signal slave_write : IN STD_LOGIC;
                    signal slave_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal master_address : OUT STD_LOGIC_VECTOR (6 DOWNTO 0);
                    signal master_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal master_nativeaddress : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
                    signal master_read : OUT STD_LOGIC;
                    signal master_write : OUT STD_LOGIC;
                    signal master_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal slave_endofpacket : OUT STD_LOGIC;
                    signal slave_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal slave_readdatavalid : OUT STD_LOGIC;
                    signal slave_waitrequest : OUT STD_LOGIC
                 );
end component clock_crossing_0;

component clock_crossing_0_bridge_arbitrator is 
end component clock_crossing_0_bridge_arbitrator;

component clock_crossing_1_s1_arbitrator is 
           port (
                 -- inputs:
                    signal ap_cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (25 DOWNTO 0);
                    signal ap_cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal ap_cpu_data_master_read : IN STD_LOGIC;
                    signal ap_cpu_data_master_waitrequest : IN STD_LOGIC;
                    signal ap_cpu_data_master_write : IN STD_LOGIC;
                    signal ap_cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal clk : IN STD_LOGIC;
                    signal clock_crossing_1_s1_endofpacket : IN STD_LOGIC;
                    signal clock_crossing_1_s1_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal clock_crossing_1_s1_readdatavalid : IN STD_LOGIC;
                    signal clock_crossing_1_s1_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal ap_cpu_data_master_granted_clock_crossing_1_s1 : OUT STD_LOGIC;
                    signal ap_cpu_data_master_qualified_request_clock_crossing_1_s1 : OUT STD_LOGIC;
                    signal ap_cpu_data_master_read_data_valid_clock_crossing_1_s1 : OUT STD_LOGIC;
                    signal ap_cpu_data_master_read_data_valid_clock_crossing_1_s1_shift_register : OUT STD_LOGIC;
                    signal ap_cpu_data_master_requests_clock_crossing_1_s1 : OUT STD_LOGIC;
                    signal clock_crossing_1_s1_address : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
                    signal clock_crossing_1_s1_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal clock_crossing_1_s1_endofpacket_from_sa : OUT STD_LOGIC;
                    signal clock_crossing_1_s1_nativeaddress : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
                    signal clock_crossing_1_s1_read : OUT STD_LOGIC;
                    signal clock_crossing_1_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal clock_crossing_1_s1_reset_n : OUT STD_LOGIC;
                    signal clock_crossing_1_s1_waitrequest_from_sa : OUT STD_LOGIC;
                    signal clock_crossing_1_s1_write : OUT STD_LOGIC;
                    signal clock_crossing_1_s1_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal d1_clock_crossing_1_s1_end_xfer : OUT STD_LOGIC
                 );
end component clock_crossing_1_s1_arbitrator;

component clock_crossing_1_m1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal clock_crossing_1_m1_address : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal clock_crossing_1_m1_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal clock_crossing_1_m1_granted_digio_pio_s1 : IN STD_LOGIC;
                    signal clock_crossing_1_m1_granted_node_switch_pio_s1 : IN STD_LOGIC;
                    signal clock_crossing_1_m1_granted_portconf_pio_s1 : IN STD_LOGIC;
                    signal clock_crossing_1_m1_granted_sync_irq_s1 : IN STD_LOGIC;
                    signal clock_crossing_1_m1_granted_sysid_control_slave : IN STD_LOGIC;
                    signal clock_crossing_1_m1_granted_system_timer_ap_s1 : IN STD_LOGIC;
                    signal clock_crossing_1_m1_qualified_request_digio_pio_s1 : IN STD_LOGIC;
                    signal clock_crossing_1_m1_qualified_request_node_switch_pio_s1 : IN STD_LOGIC;
                    signal clock_crossing_1_m1_qualified_request_portconf_pio_s1 : IN STD_LOGIC;
                    signal clock_crossing_1_m1_qualified_request_sync_irq_s1 : IN STD_LOGIC;
                    signal clock_crossing_1_m1_qualified_request_sysid_control_slave : IN STD_LOGIC;
                    signal clock_crossing_1_m1_qualified_request_system_timer_ap_s1 : IN STD_LOGIC;
                    signal clock_crossing_1_m1_read : IN STD_LOGIC;
                    signal clock_crossing_1_m1_read_data_valid_digio_pio_s1 : IN STD_LOGIC;
                    signal clock_crossing_1_m1_read_data_valid_node_switch_pio_s1 : IN STD_LOGIC;
                    signal clock_crossing_1_m1_read_data_valid_portconf_pio_s1 : IN STD_LOGIC;
                    signal clock_crossing_1_m1_read_data_valid_sync_irq_s1 : IN STD_LOGIC;
                    signal clock_crossing_1_m1_read_data_valid_sysid_control_slave : IN STD_LOGIC;
                    signal clock_crossing_1_m1_read_data_valid_system_timer_ap_s1 : IN STD_LOGIC;
                    signal clock_crossing_1_m1_requests_digio_pio_s1 : IN STD_LOGIC;
                    signal clock_crossing_1_m1_requests_node_switch_pio_s1 : IN STD_LOGIC;
                    signal clock_crossing_1_m1_requests_portconf_pio_s1 : IN STD_LOGIC;
                    signal clock_crossing_1_m1_requests_sync_irq_s1 : IN STD_LOGIC;
                    signal clock_crossing_1_m1_requests_sysid_control_slave : IN STD_LOGIC;
                    signal clock_crossing_1_m1_requests_system_timer_ap_s1 : IN STD_LOGIC;
                    signal clock_crossing_1_m1_write : IN STD_LOGIC;
                    signal clock_crossing_1_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal d1_digio_pio_s1_end_xfer : IN STD_LOGIC;
                    signal d1_node_switch_pio_s1_end_xfer : IN STD_LOGIC;
                    signal d1_portconf_pio_s1_end_xfer : IN STD_LOGIC;
                    signal d1_sync_irq_s1_end_xfer : IN STD_LOGIC;
                    signal d1_sysid_control_slave_end_xfer : IN STD_LOGIC;
                    signal d1_system_timer_ap_s1_end_xfer : IN STD_LOGIC;
                    signal digio_pio_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal node_switch_pio_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal portconf_pio_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;
                    signal sync_irq_s1_readdata_from_sa : IN STD_LOGIC;
                    signal sysid_control_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal system_timer_ap_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

                 -- outputs:
                    signal clock_crossing_1_m1_address_to_slave : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal clock_crossing_1_m1_latency_counter : OUT STD_LOGIC;
                    signal clock_crossing_1_m1_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal clock_crossing_1_m1_readdatavalid : OUT STD_LOGIC;
                    signal clock_crossing_1_m1_reset_n : OUT STD_LOGIC;
                    signal clock_crossing_1_m1_waitrequest : OUT STD_LOGIC
                 );
end component clock_crossing_1_m1_arbitrator;

component clock_crossing_1 is 
           port (
                 -- inputs:
                    signal master_clk : IN STD_LOGIC;
                    signal master_endofpacket : IN STD_LOGIC;
                    signal master_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal master_readdatavalid : IN STD_LOGIC;
                    signal master_reset_n : IN STD_LOGIC;
                    signal master_waitrequest : IN STD_LOGIC;
                    signal slave_address : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
                    signal slave_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal slave_clk : IN STD_LOGIC;
                    signal slave_nativeaddress : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
                    signal slave_read : IN STD_LOGIC;
                    signal slave_reset_n : IN STD_LOGIC;
                    signal slave_write : IN STD_LOGIC;
                    signal slave_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal master_address : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal master_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal master_nativeaddress : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
                    signal master_read : OUT STD_LOGIC;
                    signal master_write : OUT STD_LOGIC;
                    signal master_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal slave_endofpacket : OUT STD_LOGIC;
                    signal slave_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal slave_readdatavalid : OUT STD_LOGIC;
                    signal slave_waitrequest : OUT STD_LOGIC
                 );
end component clock_crossing_1;

component clock_crossing_1_bridge_arbitrator is 
end component clock_crossing_1_bridge_arbitrator;

component cnApi_Av2Av_0_ap_arbitrator is 
           port (
                 -- inputs:
                    signal ap_cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (25 DOWNTO 0);
                    signal ap_cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal ap_cpu_data_master_read : IN STD_LOGIC;
                    signal ap_cpu_data_master_waitrequest : IN STD_LOGIC;
                    signal ap_cpu_data_master_write : IN STD_LOGIC;
                    signal ap_cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal clk : IN STD_LOGIC;
                    signal cnApi_Av2Av_0_ap_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal ap_cpu_data_master_granted_cnApi_Av2Av_0_ap : OUT STD_LOGIC;
                    signal ap_cpu_data_master_qualified_request_cnApi_Av2Av_0_ap : OUT STD_LOGIC;
                    signal ap_cpu_data_master_read_data_valid_cnApi_Av2Av_0_ap : OUT STD_LOGIC;
                    signal ap_cpu_data_master_requests_cnApi_Av2Av_0_ap : OUT STD_LOGIC;
                    signal cnApi_Av2Av_0_ap_address : OUT STD_LOGIC_VECTOR (14 DOWNTO 0);
                    signal cnApi_Av2Av_0_ap_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cnApi_Av2Av_0_ap_chipselect : OUT STD_LOGIC;
                    signal cnApi_Av2Av_0_ap_read : OUT STD_LOGIC;
                    signal cnApi_Av2Av_0_ap_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal cnApi_Av2Av_0_ap_reset : OUT STD_LOGIC;
                    signal cnApi_Av2Av_0_ap_wait_counter_eq_0 : OUT STD_LOGIC;
                    signal cnApi_Av2Av_0_ap_write : OUT STD_LOGIC;
                    signal cnApi_Av2Av_0_ap_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal d1_cnApi_Av2Av_0_ap_end_xfer : OUT STD_LOGIC
                 );
end component cnApi_Av2Av_0_ap_arbitrator;

component cnApi_Av2Av_0_pcp_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cnApi_Av2Av_0_pcp_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal pcp_cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (25 DOWNTO 0);
                    signal pcp_cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal pcp_cpu_data_master_read : IN STD_LOGIC;
                    signal pcp_cpu_data_master_waitrequest : IN STD_LOGIC;
                    signal pcp_cpu_data_master_write : IN STD_LOGIC;
                    signal pcp_cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cnApi_Av2Av_0_pcp_address : OUT STD_LOGIC_VECTOR (14 DOWNTO 0);
                    signal cnApi_Av2Av_0_pcp_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cnApi_Av2Av_0_pcp_chipselect : OUT STD_LOGIC;
                    signal cnApi_Av2Av_0_pcp_read : OUT STD_LOGIC;
                    signal cnApi_Av2Av_0_pcp_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal cnApi_Av2Av_0_pcp_reset : OUT STD_LOGIC;
                    signal cnApi_Av2Av_0_pcp_wait_counter_eq_0 : OUT STD_LOGIC;
                    signal cnApi_Av2Av_0_pcp_write : OUT STD_LOGIC;
                    signal cnApi_Av2Av_0_pcp_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal d1_cnApi_Av2Av_0_pcp_end_xfer : OUT STD_LOGIC;
                    signal pcp_cpu_data_master_granted_cnApi_Av2Av_0_pcp : OUT STD_LOGIC;
                    signal pcp_cpu_data_master_qualified_request_cnApi_Av2Av_0_pcp : OUT STD_LOGIC;
                    signal pcp_cpu_data_master_read_data_valid_cnApi_Av2Av_0_pcp : OUT STD_LOGIC;
                    signal pcp_cpu_data_master_requests_cnApi_Av2Av_0_pcp : OUT STD_LOGIC
                 );
end component cnApi_Av2Av_0_pcp_arbitrator;

component cnApi_Av2Av_0 is 
           port (
                 -- inputs:
                    signal ap_Clk : IN STD_LOGIC;
                    signal ap_Reset : IN STD_LOGIC;
                    signal ap_address : IN STD_LOGIC_VECTOR (14 DOWNTO 0);
                    signal ap_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal ap_chipselect : IN STD_LOGIC;
                    signal ap_read : IN STD_LOGIC;
                    signal ap_write : IN STD_LOGIC;
                    signal ap_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal pcp_Clk : IN STD_LOGIC;
                    signal pcp_Reset : IN STD_LOGIC;
                    signal pcp_address : IN STD_LOGIC_VECTOR (14 DOWNTO 0);
                    signal pcp_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal pcp_chipselect : IN STD_LOGIC;
                    signal pcp_read : IN STD_LOGIC;
                    signal pcp_write : IN STD_LOGIC;
                    signal pcp_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal ap_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal pcp_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
                 );
end component cnApi_Av2Av_0;

component digio_pio_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal clock_crossing_1_m1_address_to_slave : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal clock_crossing_1_m1_latency_counter : IN STD_LOGIC;
                    signal clock_crossing_1_m1_nativeaddress : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
                    signal clock_crossing_1_m1_read : IN STD_LOGIC;
                    signal clock_crossing_1_m1_write : IN STD_LOGIC;
                    signal clock_crossing_1_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal digio_pio_s1_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal clock_crossing_1_m1_granted_digio_pio_s1 : OUT STD_LOGIC;
                    signal clock_crossing_1_m1_qualified_request_digio_pio_s1 : OUT STD_LOGIC;
                    signal clock_crossing_1_m1_read_data_valid_digio_pio_s1 : OUT STD_LOGIC;
                    signal clock_crossing_1_m1_requests_digio_pio_s1 : OUT STD_LOGIC;
                    signal d1_digio_pio_s1_end_xfer : OUT STD_LOGIC;
                    signal digio_pio_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal digio_pio_s1_chipselect : OUT STD_LOGIC;
                    signal digio_pio_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal digio_pio_s1_reset_n : OUT STD_LOGIC;
                    signal digio_pio_s1_write_n : OUT STD_LOGIC;
                    signal digio_pio_s1_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
                 );
end component digio_pio_s1_arbitrator;

component digio_pio is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal chipselect : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal write_n : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal bidir_port : INOUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
                 );
end component digio_pio;

component epcs_flash_controller_0_epcs_control_port_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal epcs_flash_controller_0_epcs_control_port_dataavailable : IN STD_LOGIC;
                    signal epcs_flash_controller_0_epcs_control_port_endofpacket : IN STD_LOGIC;
                    signal epcs_flash_controller_0_epcs_control_port_irq : IN STD_LOGIC;
                    signal epcs_flash_controller_0_epcs_control_port_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal epcs_flash_controller_0_epcs_control_port_readyfordata : IN STD_LOGIC;
                    signal pcp_cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (25 DOWNTO 0);
                    signal pcp_cpu_data_master_read : IN STD_LOGIC;
                    signal pcp_cpu_data_master_write : IN STD_LOGIC;
                    signal pcp_cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal pcp_cpu_instruction_master_address_to_slave : IN STD_LOGIC_VECTOR (25 DOWNTO 0);
                    signal pcp_cpu_instruction_master_latency_counter : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal pcp_cpu_instruction_master_read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal d1_epcs_flash_controller_0_epcs_control_port_end_xfer : OUT STD_LOGIC;
                    signal epcs_flash_controller_0_epcs_control_port_address : OUT STD_LOGIC_VECTOR (8 DOWNTO 0);
                    signal epcs_flash_controller_0_epcs_control_port_chipselect : OUT STD_LOGIC;
                    signal epcs_flash_controller_0_epcs_control_port_dataavailable_from_sa : OUT STD_LOGIC;
                    signal epcs_flash_controller_0_epcs_control_port_endofpacket_from_sa : OUT STD_LOGIC;
                    signal epcs_flash_controller_0_epcs_control_port_irq_from_sa : OUT STD_LOGIC;
                    signal epcs_flash_controller_0_epcs_control_port_read_n : OUT STD_LOGIC;
                    signal epcs_flash_controller_0_epcs_control_port_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal epcs_flash_controller_0_epcs_control_port_readyfordata_from_sa : OUT STD_LOGIC;
                    signal epcs_flash_controller_0_epcs_control_port_reset_n : OUT STD_LOGIC;
                    signal epcs_flash_controller_0_epcs_control_port_write_n : OUT STD_LOGIC;
                    signal epcs_flash_controller_0_epcs_control_port_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal pcp_cpu_data_master_granted_epcs_flash_controller_0_epcs_control_port : OUT STD_LOGIC;
                    signal pcp_cpu_data_master_qualified_request_epcs_flash_controller_0_epcs_control_port : OUT STD_LOGIC;
                    signal pcp_cpu_data_master_read_data_valid_epcs_flash_controller_0_epcs_control_port : OUT STD_LOGIC;
                    signal pcp_cpu_data_master_requests_epcs_flash_controller_0_epcs_control_port : OUT STD_LOGIC;
                    signal pcp_cpu_instruction_master_granted_epcs_flash_controller_0_epcs_control_port : OUT STD_LOGIC;
                    signal pcp_cpu_instruction_master_qualified_request_epcs_flash_controller_0_epcs_control_port : OUT STD_LOGIC;
                    signal pcp_cpu_instruction_master_read_data_valid_epcs_flash_controller_0_epcs_control_port : OUT STD_LOGIC;
                    signal pcp_cpu_instruction_master_requests_epcs_flash_controller_0_epcs_control_port : OUT STD_LOGIC
                 );
end component epcs_flash_controller_0_epcs_control_port_arbitrator;

component epcs_flash_controller_0 is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (8 DOWNTO 0);
                    signal chipselect : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data0 : IN STD_LOGIC;
                    signal read_n : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal write_n : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal dataavailable : OUT STD_LOGIC;
                    signal dclk : OUT STD_LOGIC;
                    signal endofpacket : OUT STD_LOGIC;
                    signal irq : OUT STD_LOGIC;
                    signal readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal readyfordata : OUT STD_LOGIC;
                    signal sce : OUT STD_LOGIC;
                    signal sdo : OUT STD_LOGIC
                 );
end component epcs_flash_controller_0;

component irq_gen_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal clock_crossing_0_m1_address_to_slave : IN STD_LOGIC_VECTOR (6 DOWNTO 0);
                    signal clock_crossing_0_m1_latency_counter : IN STD_LOGIC;
                    signal clock_crossing_0_m1_nativeaddress : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
                    signal clock_crossing_0_m1_read : IN STD_LOGIC;
                    signal clock_crossing_0_m1_write : IN STD_LOGIC;
                    signal clock_crossing_0_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal irq_gen_s1_readdata : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal clock_crossing_0_m1_granted_irq_gen_s1 : OUT STD_LOGIC;
                    signal clock_crossing_0_m1_qualified_request_irq_gen_s1 : OUT STD_LOGIC;
                    signal clock_crossing_0_m1_read_data_valid_irq_gen_s1 : OUT STD_LOGIC;
                    signal clock_crossing_0_m1_requests_irq_gen_s1 : OUT STD_LOGIC;
                    signal d1_irq_gen_s1_end_xfer : OUT STD_LOGIC;
                    signal irq_gen_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal irq_gen_s1_chipselect : OUT STD_LOGIC;
                    signal irq_gen_s1_readdata_from_sa : OUT STD_LOGIC;
                    signal irq_gen_s1_reset_n : OUT STD_LOGIC;
                    signal irq_gen_s1_write_n : OUT STD_LOGIC;
                    signal irq_gen_s1_writedata : OUT STD_LOGIC
                 );
end component irq_gen_s1_arbitrator;

component irq_gen is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal chipselect : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal write_n : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC;

                 -- outputs:
                    signal out_port : OUT STD_LOGIC;
                    signal readdata : OUT STD_LOGIC
                 );
end component irq_gen;

component jtag_uart_0_avalon_jtag_slave_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal jtag_uart_0_avalon_jtag_slave_dataavailable : IN STD_LOGIC;
                    signal jtag_uart_0_avalon_jtag_slave_irq : IN STD_LOGIC;
                    signal jtag_uart_0_avalon_jtag_slave_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal jtag_uart_0_avalon_jtag_slave_readyfordata : IN STD_LOGIC;
                    signal jtag_uart_0_avalon_jtag_slave_waitrequest : IN STD_LOGIC;
                    signal niosII_openMac_clock_0_out_address_to_slave : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal niosII_openMac_clock_0_out_nativeaddress : IN STD_LOGIC;
                    signal niosII_openMac_clock_0_out_read : IN STD_LOGIC;
                    signal niosII_openMac_clock_0_out_write : IN STD_LOGIC;
                    signal niosII_openMac_clock_0_out_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal d1_jtag_uart_0_avalon_jtag_slave_end_xfer : OUT STD_LOGIC;
                    signal jtag_uart_0_avalon_jtag_slave_address : OUT STD_LOGIC;
                    signal jtag_uart_0_avalon_jtag_slave_chipselect : OUT STD_LOGIC;
                    signal jtag_uart_0_avalon_jtag_slave_dataavailable_from_sa : OUT STD_LOGIC;
                    signal jtag_uart_0_avalon_jtag_slave_irq_from_sa : OUT STD_LOGIC;
                    signal jtag_uart_0_avalon_jtag_slave_read_n : OUT STD_LOGIC;
                    signal jtag_uart_0_avalon_jtag_slave_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal jtag_uart_0_avalon_jtag_slave_readyfordata_from_sa : OUT STD_LOGIC;
                    signal jtag_uart_0_avalon_jtag_slave_reset_n : OUT STD_LOGIC;
                    signal jtag_uart_0_avalon_jtag_slave_waitrequest_from_sa : OUT STD_LOGIC;
                    signal jtag_uart_0_avalon_jtag_slave_write_n : OUT STD_LOGIC;
                    signal jtag_uart_0_avalon_jtag_slave_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal niosII_openMac_clock_0_out_granted_jtag_uart_0_avalon_jtag_slave : OUT STD_LOGIC;
                    signal niosII_openMac_clock_0_out_qualified_request_jtag_uart_0_avalon_jtag_slave : OUT STD_LOGIC;
                    signal niosII_openMac_clock_0_out_read_data_valid_jtag_uart_0_avalon_jtag_slave : OUT STD_LOGIC;
                    signal niosII_openMac_clock_0_out_requests_jtag_uart_0_avalon_jtag_slave : OUT STD_LOGIC
                 );
end component jtag_uart_0_avalon_jtag_slave_arbitrator;

component jtag_uart_0 is 
           port (
                 -- inputs:
                    signal av_address : IN STD_LOGIC;
                    signal av_chipselect : IN STD_LOGIC;
                    signal av_read_n : IN STD_LOGIC;
                    signal av_write_n : IN STD_LOGIC;
                    signal av_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal clk : IN STD_LOGIC;
                    signal rst_n : IN STD_LOGIC;

                 -- outputs:
                    signal av_irq : OUT STD_LOGIC;
                    signal av_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal av_waitrequest : OUT STD_LOGIC;
                    signal dataavailable : OUT STD_LOGIC;
                    signal readyfordata : OUT STD_LOGIC
                 );
end component jtag_uart_0;

component jtag_uart_1_avalon_jtag_slave_arbitrator is 
           port (
                 -- inputs:
                    signal ap_cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (25 DOWNTO 0);
                    signal ap_cpu_data_master_read : IN STD_LOGIC;
                    signal ap_cpu_data_master_waitrequest : IN STD_LOGIC;
                    signal ap_cpu_data_master_write : IN STD_LOGIC;
                    signal ap_cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal clk : IN STD_LOGIC;
                    signal jtag_uart_1_avalon_jtag_slave_dataavailable : IN STD_LOGIC;
                    signal jtag_uart_1_avalon_jtag_slave_irq : IN STD_LOGIC;
                    signal jtag_uart_1_avalon_jtag_slave_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal jtag_uart_1_avalon_jtag_slave_readyfordata : IN STD_LOGIC;
                    signal jtag_uart_1_avalon_jtag_slave_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal ap_cpu_data_master_granted_jtag_uart_1_avalon_jtag_slave : OUT STD_LOGIC;
                    signal ap_cpu_data_master_qualified_request_jtag_uart_1_avalon_jtag_slave : OUT STD_LOGIC;
                    signal ap_cpu_data_master_read_data_valid_jtag_uart_1_avalon_jtag_slave : OUT STD_LOGIC;
                    signal ap_cpu_data_master_requests_jtag_uart_1_avalon_jtag_slave : OUT STD_LOGIC;
                    signal d1_jtag_uart_1_avalon_jtag_slave_end_xfer : OUT STD_LOGIC;
                    signal jtag_uart_1_avalon_jtag_slave_address : OUT STD_LOGIC;
                    signal jtag_uart_1_avalon_jtag_slave_chipselect : OUT STD_LOGIC;
                    signal jtag_uart_1_avalon_jtag_slave_dataavailable_from_sa : OUT STD_LOGIC;
                    signal jtag_uart_1_avalon_jtag_slave_irq_from_sa : OUT STD_LOGIC;
                    signal jtag_uart_1_avalon_jtag_slave_read_n : OUT STD_LOGIC;
                    signal jtag_uart_1_avalon_jtag_slave_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal jtag_uart_1_avalon_jtag_slave_readyfordata_from_sa : OUT STD_LOGIC;
                    signal jtag_uart_1_avalon_jtag_slave_reset_n : OUT STD_LOGIC;
                    signal jtag_uart_1_avalon_jtag_slave_waitrequest_from_sa : OUT STD_LOGIC;
                    signal jtag_uart_1_avalon_jtag_slave_write_n : OUT STD_LOGIC;
                    signal jtag_uart_1_avalon_jtag_slave_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
                 );
end component jtag_uart_1_avalon_jtag_slave_arbitrator;

component jtag_uart_1 is 
           port (
                 -- inputs:
                    signal av_address : IN STD_LOGIC;
                    signal av_chipselect : IN STD_LOGIC;
                    signal av_read_n : IN STD_LOGIC;
                    signal av_write_n : IN STD_LOGIC;
                    signal av_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal clk : IN STD_LOGIC;
                    signal rst_n : IN STD_LOGIC;

                 -- outputs:
                    signal av_irq : OUT STD_LOGIC;
                    signal av_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal av_waitrequest : OUT STD_LOGIC;
                    signal dataavailable : OUT STD_LOGIC;
                    signal readyfordata : OUT STD_LOGIC
                 );
end component jtag_uart_1;

component niosII_openMac_clock_0_in_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal niosII_openMac_clock_0_in_endofpacket : IN STD_LOGIC;
                    signal niosII_openMac_clock_0_in_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal niosII_openMac_clock_0_in_waitrequest : IN STD_LOGIC;
                    signal pcp_cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (25 DOWNTO 0);
                    signal pcp_cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal pcp_cpu_data_master_read : IN STD_LOGIC;
                    signal pcp_cpu_data_master_waitrequest : IN STD_LOGIC;
                    signal pcp_cpu_data_master_write : IN STD_LOGIC;
                    signal pcp_cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal d1_niosII_openMac_clock_0_in_end_xfer : OUT STD_LOGIC;
                    signal niosII_openMac_clock_0_in_address : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal niosII_openMac_clock_0_in_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal niosII_openMac_clock_0_in_endofpacket_from_sa : OUT STD_LOGIC;
                    signal niosII_openMac_clock_0_in_nativeaddress : OUT STD_LOGIC;
                    signal niosII_openMac_clock_0_in_read : OUT STD_LOGIC;
                    signal niosII_openMac_clock_0_in_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal niosII_openMac_clock_0_in_reset_n : OUT STD_LOGIC;
                    signal niosII_openMac_clock_0_in_waitrequest_from_sa : OUT STD_LOGIC;
                    signal niosII_openMac_clock_0_in_write : OUT STD_LOGIC;
                    signal niosII_openMac_clock_0_in_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal pcp_cpu_data_master_granted_niosII_openMac_clock_0_in : OUT STD_LOGIC;
                    signal pcp_cpu_data_master_qualified_request_niosII_openMac_clock_0_in : OUT STD_LOGIC;
                    signal pcp_cpu_data_master_read_data_valid_niosII_openMac_clock_0_in : OUT STD_LOGIC;
                    signal pcp_cpu_data_master_requests_niosII_openMac_clock_0_in : OUT STD_LOGIC
                 );
end component niosII_openMac_clock_0_in_arbitrator;

component niosII_openMac_clock_0_out_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal d1_jtag_uart_0_avalon_jtag_slave_end_xfer : IN STD_LOGIC;
                    signal jtag_uart_0_avalon_jtag_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal jtag_uart_0_avalon_jtag_slave_waitrequest_from_sa : IN STD_LOGIC;
                    signal niosII_openMac_clock_0_out_address : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal niosII_openMac_clock_0_out_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal niosII_openMac_clock_0_out_granted_jtag_uart_0_avalon_jtag_slave : IN STD_LOGIC;
                    signal niosII_openMac_clock_0_out_qualified_request_jtag_uart_0_avalon_jtag_slave : IN STD_LOGIC;
                    signal niosII_openMac_clock_0_out_read : IN STD_LOGIC;
                    signal niosII_openMac_clock_0_out_read_data_valid_jtag_uart_0_avalon_jtag_slave : IN STD_LOGIC;
                    signal niosII_openMac_clock_0_out_requests_jtag_uart_0_avalon_jtag_slave : IN STD_LOGIC;
                    signal niosII_openMac_clock_0_out_write : IN STD_LOGIC;
                    signal niosII_openMac_clock_0_out_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal niosII_openMac_clock_0_out_address_to_slave : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal niosII_openMac_clock_0_out_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal niosII_openMac_clock_0_out_reset_n : OUT STD_LOGIC;
                    signal niosII_openMac_clock_0_out_waitrequest : OUT STD_LOGIC
                 );
end component niosII_openMac_clock_0_out_arbitrator;

component niosII_openMac_clock_0 is 
           port (
                 -- inputs:
                    signal master_clk : IN STD_LOGIC;
                    signal master_endofpacket : IN STD_LOGIC;
                    signal master_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal master_reset_n : IN STD_LOGIC;
                    signal master_waitrequest : IN STD_LOGIC;
                    signal slave_address : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal slave_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal slave_clk : IN STD_LOGIC;
                    signal slave_nativeaddress : IN STD_LOGIC;
                    signal slave_read : IN STD_LOGIC;
                    signal slave_reset_n : IN STD_LOGIC;
                    signal slave_write : IN STD_LOGIC;
                    signal slave_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal master_address : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal master_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal master_nativeaddress : OUT STD_LOGIC;
                    signal master_read : OUT STD_LOGIC;
                    signal master_write : OUT STD_LOGIC;
                    signal master_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal slave_endofpacket : OUT STD_LOGIC;
                    signal slave_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal slave_waitrequest : OUT STD_LOGIC
                 );
end component niosII_openMac_clock_0;

component niosII_openMac_clock_1_in_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal niosII_openMac_clock_1_in_endofpacket : IN STD_LOGIC;
                    signal niosII_openMac_clock_1_in_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal niosII_openMac_clock_1_in_waitrequest : IN STD_LOGIC;
                    signal pcp_cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (25 DOWNTO 0);
                    signal pcp_cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal pcp_cpu_data_master_read : IN STD_LOGIC;
                    signal pcp_cpu_data_master_waitrequest : IN STD_LOGIC;
                    signal pcp_cpu_data_master_write : IN STD_LOGIC;
                    signal pcp_cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal d1_niosII_openMac_clock_1_in_end_xfer : OUT STD_LOGIC;
                    signal niosII_openMac_clock_1_in_address : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal niosII_openMac_clock_1_in_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal niosII_openMac_clock_1_in_endofpacket_from_sa : OUT STD_LOGIC;
                    signal niosII_openMac_clock_1_in_nativeaddress : OUT STD_LOGIC;
                    signal niosII_openMac_clock_1_in_read : OUT STD_LOGIC;
                    signal niosII_openMac_clock_1_in_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal niosII_openMac_clock_1_in_reset_n : OUT STD_LOGIC;
                    signal niosII_openMac_clock_1_in_waitrequest_from_sa : OUT STD_LOGIC;
                    signal niosII_openMac_clock_1_in_write : OUT STD_LOGIC;
                    signal niosII_openMac_clock_1_in_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal pcp_cpu_data_master_granted_niosII_openMac_clock_1_in : OUT STD_LOGIC;
                    signal pcp_cpu_data_master_qualified_request_niosII_openMac_clock_1_in : OUT STD_LOGIC;
                    signal pcp_cpu_data_master_read_data_valid_niosII_openMac_clock_1_in : OUT STD_LOGIC;
                    signal pcp_cpu_data_master_requests_niosII_openMac_clock_1_in : OUT STD_LOGIC
                 );
end component niosII_openMac_clock_1_in_arbitrator;

component niosII_openMac_clock_1_out_arbitrator is 
           port (
                 -- inputs:
                    signal OpenMAC_0_CMP_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal clk : IN STD_LOGIC;
                    signal d1_OpenMAC_0_CMP_end_xfer : IN STD_LOGIC;
                    signal niosII_openMac_clock_1_out_address : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal niosII_openMac_clock_1_out_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal niosII_openMac_clock_1_out_granted_OpenMAC_0_CMP : IN STD_LOGIC;
                    signal niosII_openMac_clock_1_out_qualified_request_OpenMAC_0_CMP : IN STD_LOGIC;
                    signal niosII_openMac_clock_1_out_read : IN STD_LOGIC;
                    signal niosII_openMac_clock_1_out_read_data_valid_OpenMAC_0_CMP : IN STD_LOGIC;
                    signal niosII_openMac_clock_1_out_requests_OpenMAC_0_CMP : IN STD_LOGIC;
                    signal niosII_openMac_clock_1_out_write : IN STD_LOGIC;
                    signal niosII_openMac_clock_1_out_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal niosII_openMac_clock_1_out_address_to_slave : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal niosII_openMac_clock_1_out_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal niosII_openMac_clock_1_out_reset_n : OUT STD_LOGIC;
                    signal niosII_openMac_clock_1_out_waitrequest : OUT STD_LOGIC
                 );
end component niosII_openMac_clock_1_out_arbitrator;

component niosII_openMac_clock_1 is 
           port (
                 -- inputs:
                    signal master_clk : IN STD_LOGIC;
                    signal master_endofpacket : IN STD_LOGIC;
                    signal master_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal master_reset_n : IN STD_LOGIC;
                    signal master_waitrequest : IN STD_LOGIC;
                    signal slave_address : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal slave_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal slave_clk : IN STD_LOGIC;
                    signal slave_nativeaddress : IN STD_LOGIC;
                    signal slave_read : IN STD_LOGIC;
                    signal slave_reset_n : IN STD_LOGIC;
                    signal slave_write : IN STD_LOGIC;
                    signal slave_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal master_address : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal master_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal master_nativeaddress : OUT STD_LOGIC;
                    signal master_read : OUT STD_LOGIC;
                    signal master_write : OUT STD_LOGIC;
                    signal master_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal slave_endofpacket : OUT STD_LOGIC;
                    signal slave_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal slave_waitrequest : OUT STD_LOGIC
                 );
end component niosII_openMac_clock_1;

component niosII_openMac_clock_2_in_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal niosII_openMac_clock_2_in_endofpacket : IN STD_LOGIC;
                    signal niosII_openMac_clock_2_in_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal niosII_openMac_clock_2_in_waitrequest : IN STD_LOGIC;
                    signal pcp_cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (25 DOWNTO 0);
                    signal pcp_cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal pcp_cpu_data_master_dbs_address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal pcp_cpu_data_master_dbs_write_16 : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal pcp_cpu_data_master_no_byte_enables_and_last_term : IN STD_LOGIC;
                    signal pcp_cpu_data_master_read : IN STD_LOGIC;
                    signal pcp_cpu_data_master_waitrequest : IN STD_LOGIC;
                    signal pcp_cpu_data_master_write : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal d1_niosII_openMac_clock_2_in_end_xfer : OUT STD_LOGIC;
                    signal niosII_openMac_clock_2_in_address : OUT STD_LOGIC_VECTOR (12 DOWNTO 0);
                    signal niosII_openMac_clock_2_in_byteenable : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal niosII_openMac_clock_2_in_endofpacket_from_sa : OUT STD_LOGIC;
                    signal niosII_openMac_clock_2_in_nativeaddress : OUT STD_LOGIC_VECTOR (11 DOWNTO 0);
                    signal niosII_openMac_clock_2_in_read : OUT STD_LOGIC;
                    signal niosII_openMac_clock_2_in_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal niosII_openMac_clock_2_in_reset_n : OUT STD_LOGIC;
                    signal niosII_openMac_clock_2_in_waitrequest_from_sa : OUT STD_LOGIC;
                    signal niosII_openMac_clock_2_in_write : OUT STD_LOGIC;
                    signal niosII_openMac_clock_2_in_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal pcp_cpu_data_master_byteenable_niosII_openMac_clock_2_in : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal pcp_cpu_data_master_granted_niosII_openMac_clock_2_in : OUT STD_LOGIC;
                    signal pcp_cpu_data_master_qualified_request_niosII_openMac_clock_2_in : OUT STD_LOGIC;
                    signal pcp_cpu_data_master_read_data_valid_niosII_openMac_clock_2_in : OUT STD_LOGIC;
                    signal pcp_cpu_data_master_requests_niosII_openMac_clock_2_in : OUT STD_LOGIC
                 );
end component niosII_openMac_clock_2_in_arbitrator;

component niosII_openMac_clock_2_out_arbitrator is 
           port (
                 -- inputs:
                    signal OpenMAC_0_REG_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal clk : IN STD_LOGIC;
                    signal d1_OpenMAC_0_REG_end_xfer : IN STD_LOGIC;
                    signal niosII_openMac_clock_2_out_address : IN STD_LOGIC_VECTOR (12 DOWNTO 0);
                    signal niosII_openMac_clock_2_out_byteenable : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal niosII_openMac_clock_2_out_granted_OpenMAC_0_REG : IN STD_LOGIC;
                    signal niosII_openMac_clock_2_out_qualified_request_OpenMAC_0_REG : IN STD_LOGIC;
                    signal niosII_openMac_clock_2_out_read : IN STD_LOGIC;
                    signal niosII_openMac_clock_2_out_read_data_valid_OpenMAC_0_REG : IN STD_LOGIC;
                    signal niosII_openMac_clock_2_out_requests_OpenMAC_0_REG : IN STD_LOGIC;
                    signal niosII_openMac_clock_2_out_write : IN STD_LOGIC;
                    signal niosII_openMac_clock_2_out_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal niosII_openMac_clock_2_out_address_to_slave : OUT STD_LOGIC_VECTOR (12 DOWNTO 0);
                    signal niosII_openMac_clock_2_out_readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal niosII_openMac_clock_2_out_reset_n : OUT STD_LOGIC;
                    signal niosII_openMac_clock_2_out_waitrequest : OUT STD_LOGIC
                 );
end component niosII_openMac_clock_2_out_arbitrator;

component niosII_openMac_clock_2 is 
           port (
                 -- inputs:
                    signal master_clk : IN STD_LOGIC;
                    signal master_endofpacket : IN STD_LOGIC;
                    signal master_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal master_reset_n : IN STD_LOGIC;
                    signal master_waitrequest : IN STD_LOGIC;
                    signal slave_address : IN STD_LOGIC_VECTOR (12 DOWNTO 0);
                    signal slave_byteenable : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal slave_clk : IN STD_LOGIC;
                    signal slave_nativeaddress : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
                    signal slave_read : IN STD_LOGIC;
                    signal slave_reset_n : IN STD_LOGIC;
                    signal slave_write : IN STD_LOGIC;
                    signal slave_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

                 -- outputs:
                    signal master_address : OUT STD_LOGIC_VECTOR (12 DOWNTO 0);
                    signal master_byteenable : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal master_nativeaddress : OUT STD_LOGIC_VECTOR (11 DOWNTO 0);
                    signal master_read : OUT STD_LOGIC;
                    signal master_write : OUT STD_LOGIC;
                    signal master_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal slave_endofpacket : OUT STD_LOGIC;
                    signal slave_readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal slave_waitrequest : OUT STD_LOGIC
                 );
end component niosII_openMac_clock_2;

component niosII_openMac_clock_3_in_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal niosII_openMac_clock_3_in_endofpacket : IN STD_LOGIC;
                    signal niosII_openMac_clock_3_in_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal niosII_openMac_clock_3_in_waitrequest : IN STD_LOGIC;
                    signal pcp_cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (25 DOWNTO 0);
                    signal pcp_cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal pcp_cpu_data_master_read : IN STD_LOGIC;
                    signal pcp_cpu_data_master_waitrequest : IN STD_LOGIC;
                    signal pcp_cpu_data_master_write : IN STD_LOGIC;
                    signal pcp_cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal d1_niosII_openMac_clock_3_in_end_xfer : OUT STD_LOGIC;
                    signal niosII_openMac_clock_3_in_address : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal niosII_openMac_clock_3_in_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal niosII_openMac_clock_3_in_endofpacket_from_sa : OUT STD_LOGIC;
                    signal niosII_openMac_clock_3_in_nativeaddress : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal niosII_openMac_clock_3_in_read : OUT STD_LOGIC;
                    signal niosII_openMac_clock_3_in_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal niosII_openMac_clock_3_in_reset_n : OUT STD_LOGIC;
                    signal niosII_openMac_clock_3_in_waitrequest_from_sa : OUT STD_LOGIC;
                    signal niosII_openMac_clock_3_in_write : OUT STD_LOGIC;
                    signal niosII_openMac_clock_3_in_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal pcp_cpu_data_master_granted_niosII_openMac_clock_3_in : OUT STD_LOGIC;
                    signal pcp_cpu_data_master_qualified_request_niosII_openMac_clock_3_in : OUT STD_LOGIC;
                    signal pcp_cpu_data_master_read_data_valid_niosII_openMac_clock_3_in : OUT STD_LOGIC;
                    signal pcp_cpu_data_master_requests_niosII_openMac_clock_3_in : OUT STD_LOGIC
                 );
end component niosII_openMac_clock_3_in_arbitrator;

component niosII_openMac_clock_3_out_arbitrator is 
           port (
                 -- inputs:
                    signal altpll_0_pll_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal clk : IN STD_LOGIC;
                    signal d1_altpll_0_pll_slave_end_xfer : IN STD_LOGIC;
                    signal niosII_openMac_clock_3_out_address : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal niosII_openMac_clock_3_out_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal niosII_openMac_clock_3_out_granted_altpll_0_pll_slave : IN STD_LOGIC;
                    signal niosII_openMac_clock_3_out_qualified_request_altpll_0_pll_slave : IN STD_LOGIC;
                    signal niosII_openMac_clock_3_out_read : IN STD_LOGIC;
                    signal niosII_openMac_clock_3_out_read_data_valid_altpll_0_pll_slave : IN STD_LOGIC;
                    signal niosII_openMac_clock_3_out_requests_altpll_0_pll_slave : IN STD_LOGIC;
                    signal niosII_openMac_clock_3_out_write : IN STD_LOGIC;
                    signal niosII_openMac_clock_3_out_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal niosII_openMac_clock_3_out_address_to_slave : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal niosII_openMac_clock_3_out_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal niosII_openMac_clock_3_out_reset_n : OUT STD_LOGIC;
                    signal niosII_openMac_clock_3_out_waitrequest : OUT STD_LOGIC
                 );
end component niosII_openMac_clock_3_out_arbitrator;

component niosII_openMac_clock_3 is 
           port (
                 -- inputs:
                    signal master_clk : IN STD_LOGIC;
                    signal master_endofpacket : IN STD_LOGIC;
                    signal master_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal master_reset_n : IN STD_LOGIC;
                    signal master_waitrequest : IN STD_LOGIC;
                    signal slave_address : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal slave_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal slave_clk : IN STD_LOGIC;
                    signal slave_nativeaddress : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal slave_read : IN STD_LOGIC;
                    signal slave_reset_n : IN STD_LOGIC;
                    signal slave_write : IN STD_LOGIC;
                    signal slave_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal master_address : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal master_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal master_nativeaddress : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal master_read : OUT STD_LOGIC;
                    signal master_write : OUT STD_LOGIC;
                    signal master_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal slave_endofpacket : OUT STD_LOGIC;
                    signal slave_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal slave_waitrequest : OUT STD_LOGIC
                 );
end component niosII_openMac_clock_3;

component niosII_openMac_clock_4_in_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal niosII_openMac_clock_4_in_endofpacket : IN STD_LOGIC;
                    signal niosII_openMac_clock_4_in_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal niosII_openMac_clock_4_in_waitrequest : IN STD_LOGIC;
                    signal pcp_cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (25 DOWNTO 0);
                    signal pcp_cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal pcp_cpu_data_master_read : IN STD_LOGIC;
                    signal pcp_cpu_data_master_waitrequest : IN STD_LOGIC;
                    signal pcp_cpu_data_master_write : IN STD_LOGIC;
                    signal pcp_cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal d1_niosII_openMac_clock_4_in_end_xfer : OUT STD_LOGIC;
                    signal niosII_openMac_clock_4_in_address : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal niosII_openMac_clock_4_in_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal niosII_openMac_clock_4_in_endofpacket_from_sa : OUT STD_LOGIC;
                    signal niosII_openMac_clock_4_in_nativeaddress : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
                    signal niosII_openMac_clock_4_in_read : OUT STD_LOGIC;
                    signal niosII_openMac_clock_4_in_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal niosII_openMac_clock_4_in_reset_n : OUT STD_LOGIC;
                    signal niosII_openMac_clock_4_in_waitrequest_from_sa : OUT STD_LOGIC;
                    signal niosII_openMac_clock_4_in_write : OUT STD_LOGIC;
                    signal niosII_openMac_clock_4_in_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal pcp_cpu_data_master_granted_niosII_openMac_clock_4_in : OUT STD_LOGIC;
                    signal pcp_cpu_data_master_qualified_request_niosII_openMac_clock_4_in : OUT STD_LOGIC;
                    signal pcp_cpu_data_master_read_data_valid_niosII_openMac_clock_4_in : OUT STD_LOGIC;
                    signal pcp_cpu_data_master_requests_niosII_openMac_clock_4_in : OUT STD_LOGIC
                 );
end component niosII_openMac_clock_4_in_arbitrator;

component niosII_openMac_clock_4_out_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal d1_remote_update_cycloneiii_0_s1_end_xfer : IN STD_LOGIC;
                    signal niosII_openMac_clock_4_out_address : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal niosII_openMac_clock_4_out_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal niosII_openMac_clock_4_out_granted_remote_update_cycloneiii_0_s1 : IN STD_LOGIC;
                    signal niosII_openMac_clock_4_out_qualified_request_remote_update_cycloneiii_0_s1 : IN STD_LOGIC;
                    signal niosII_openMac_clock_4_out_read : IN STD_LOGIC;
                    signal niosII_openMac_clock_4_out_read_data_valid_remote_update_cycloneiii_0_s1 : IN STD_LOGIC;
                    signal niosII_openMac_clock_4_out_requests_remote_update_cycloneiii_0_s1 : IN STD_LOGIC;
                    signal niosII_openMac_clock_4_out_write : IN STD_LOGIC;
                    signal niosII_openMac_clock_4_out_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal remote_update_cycloneiii_0_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal remote_update_cycloneiii_0_s1_waitrequest_from_sa : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal niosII_openMac_clock_4_out_address_to_slave : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal niosII_openMac_clock_4_out_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal niosII_openMac_clock_4_out_reset_n : OUT STD_LOGIC;
                    signal niosII_openMac_clock_4_out_waitrequest : OUT STD_LOGIC
                 );
end component niosII_openMac_clock_4_out_arbitrator;

component niosII_openMac_clock_4 is 
           port (
                 -- inputs:
                    signal master_clk : IN STD_LOGIC;
                    signal master_endofpacket : IN STD_LOGIC;
                    signal master_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal master_reset_n : IN STD_LOGIC;
                    signal master_waitrequest : IN STD_LOGIC;
                    signal slave_address : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal slave_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal slave_clk : IN STD_LOGIC;
                    signal slave_nativeaddress : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
                    signal slave_read : IN STD_LOGIC;
                    signal slave_reset_n : IN STD_LOGIC;
                    signal slave_write : IN STD_LOGIC;
                    signal slave_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal master_address : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal master_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal master_nativeaddress : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
                    signal master_read : OUT STD_LOGIC;
                    signal master_write : OUT STD_LOGIC;
                    signal master_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal slave_endofpacket : OUT STD_LOGIC;
                    signal slave_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal slave_waitrequest : OUT STD_LOGIC
                 );
end component niosII_openMac_clock_4;

component node_switch_pio_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal clock_crossing_1_m1_address_to_slave : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal clock_crossing_1_m1_latency_counter : IN STD_LOGIC;
                    signal clock_crossing_1_m1_nativeaddress : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
                    signal clock_crossing_1_m1_read : IN STD_LOGIC;
                    signal clock_crossing_1_m1_write : IN STD_LOGIC;
                    signal node_switch_pio_s1_readdata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal clock_crossing_1_m1_granted_node_switch_pio_s1 : OUT STD_LOGIC;
                    signal clock_crossing_1_m1_qualified_request_node_switch_pio_s1 : OUT STD_LOGIC;
                    signal clock_crossing_1_m1_read_data_valid_node_switch_pio_s1 : OUT STD_LOGIC;
                    signal clock_crossing_1_m1_requests_node_switch_pio_s1 : OUT STD_LOGIC;
                    signal d1_node_switch_pio_s1_end_xfer : OUT STD_LOGIC;
                    signal node_switch_pio_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal node_switch_pio_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal node_switch_pio_s1_reset_n : OUT STD_LOGIC
                 );
end component node_switch_pio_s1_arbitrator;

component node_switch_pio is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal clk : IN STD_LOGIC;
                    signal in_port : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal readdata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
                 );
end component node_switch_pio;

component onchip_memory_0_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal onchip_memory_0_s1_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal pcp_cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (25 DOWNTO 0);
                    signal pcp_cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal pcp_cpu_data_master_read : IN STD_LOGIC;
                    signal pcp_cpu_data_master_waitrequest : IN STD_LOGIC;
                    signal pcp_cpu_data_master_write : IN STD_LOGIC;
                    signal pcp_cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal pcp_cpu_instruction_master_address_to_slave : IN STD_LOGIC_VECTOR (25 DOWNTO 0);
                    signal pcp_cpu_instruction_master_latency_counter : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal pcp_cpu_instruction_master_read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal d1_onchip_memory_0_s1_end_xfer : OUT STD_LOGIC;
                    signal onchip_memory_0_s1_address : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal onchip_memory_0_s1_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal onchip_memory_0_s1_chipselect : OUT STD_LOGIC;
                    signal onchip_memory_0_s1_clken : OUT STD_LOGIC;
                    signal onchip_memory_0_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal onchip_memory_0_s1_write : OUT STD_LOGIC;
                    signal onchip_memory_0_s1_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal pcp_cpu_data_master_granted_onchip_memory_0_s1 : OUT STD_LOGIC;
                    signal pcp_cpu_data_master_qualified_request_onchip_memory_0_s1 : OUT STD_LOGIC;
                    signal pcp_cpu_data_master_read_data_valid_onchip_memory_0_s1 : OUT STD_LOGIC;
                    signal pcp_cpu_data_master_requests_onchip_memory_0_s1 : OUT STD_LOGIC;
                    signal pcp_cpu_instruction_master_granted_onchip_memory_0_s1 : OUT STD_LOGIC;
                    signal pcp_cpu_instruction_master_qualified_request_onchip_memory_0_s1 : OUT STD_LOGIC;
                    signal pcp_cpu_instruction_master_read_data_valid_onchip_memory_0_s1 : OUT STD_LOGIC;
                    signal pcp_cpu_instruction_master_requests_onchip_memory_0_s1 : OUT STD_LOGIC;
                    signal registered_pcp_cpu_data_master_read_data_valid_onchip_memory_0_s1 : OUT STD_LOGIC
                 );
end component onchip_memory_0_s1_arbitrator;

component onchip_memory_0 is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal chipselect : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal clken : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
                 );
end component onchip_memory_0;

component pcp_cpu_jtag_debug_module_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal pcp_cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (25 DOWNTO 0);
                    signal pcp_cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal pcp_cpu_data_master_debugaccess : IN STD_LOGIC;
                    signal pcp_cpu_data_master_read : IN STD_LOGIC;
                    signal pcp_cpu_data_master_waitrequest : IN STD_LOGIC;
                    signal pcp_cpu_data_master_write : IN STD_LOGIC;
                    signal pcp_cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal pcp_cpu_instruction_master_address_to_slave : IN STD_LOGIC_VECTOR (25 DOWNTO 0);
                    signal pcp_cpu_instruction_master_latency_counter : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal pcp_cpu_instruction_master_read : IN STD_LOGIC;
                    signal pcp_cpu_jtag_debug_module_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal pcp_cpu_jtag_debug_module_resetrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal d1_pcp_cpu_jtag_debug_module_end_xfer : OUT STD_LOGIC;
                    signal pcp_cpu_data_master_granted_pcp_cpu_jtag_debug_module : OUT STD_LOGIC;
                    signal pcp_cpu_data_master_qualified_request_pcp_cpu_jtag_debug_module : OUT STD_LOGIC;
                    signal pcp_cpu_data_master_read_data_valid_pcp_cpu_jtag_debug_module : OUT STD_LOGIC;
                    signal pcp_cpu_data_master_requests_pcp_cpu_jtag_debug_module : OUT STD_LOGIC;
                    signal pcp_cpu_instruction_master_granted_pcp_cpu_jtag_debug_module : OUT STD_LOGIC;
                    signal pcp_cpu_instruction_master_qualified_request_pcp_cpu_jtag_debug_module : OUT STD_LOGIC;
                    signal pcp_cpu_instruction_master_read_data_valid_pcp_cpu_jtag_debug_module : OUT STD_LOGIC;
                    signal pcp_cpu_instruction_master_requests_pcp_cpu_jtag_debug_module : OUT STD_LOGIC;
                    signal pcp_cpu_jtag_debug_module_address : OUT STD_LOGIC_VECTOR (8 DOWNTO 0);
                    signal pcp_cpu_jtag_debug_module_begintransfer : OUT STD_LOGIC;
                    signal pcp_cpu_jtag_debug_module_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal pcp_cpu_jtag_debug_module_chipselect : OUT STD_LOGIC;
                    signal pcp_cpu_jtag_debug_module_debugaccess : OUT STD_LOGIC;
                    signal pcp_cpu_jtag_debug_module_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal pcp_cpu_jtag_debug_module_reset_n : OUT STD_LOGIC;
                    signal pcp_cpu_jtag_debug_module_resetrequest_from_sa : OUT STD_LOGIC;
                    signal pcp_cpu_jtag_debug_module_write : OUT STD_LOGIC;
                    signal pcp_cpu_jtag_debug_module_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
                 );
end component pcp_cpu_jtag_debug_module_arbitrator;

component pcp_cpu_data_master_arbitrator is 
           port (
                 -- inputs:
                    signal DBC3C40_SRAM_0_avalon_tristate_slave_wait_counter_eq_0 : IN STD_LOGIC;
                    signal OpenMAC_0_CMP_irq_from_sa : IN STD_LOGIC;
                    signal OpenMAC_0_REG_irq_from_sa : IN STD_LOGIC;
                    signal OpenMAC_0_iBuf_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal OpenMAC_0_iBuf_wait_counter_eq_0 : IN STD_LOGIC;
                    signal cfi_flash_0_s1_wait_counter_eq_0 : IN STD_LOGIC;
                    signal cfi_flash_0_s1_wait_counter_eq_1 : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal clk90Meg : IN STD_LOGIC;
                    signal clk90Meg_reset_n : IN STD_LOGIC;
                    signal clock_crossing_0_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal clock_crossing_0_s1_waitrequest_from_sa : IN STD_LOGIC;
                    signal cnApi_Av2Av_0_pcp_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal cnApi_Av2Av_0_pcp_wait_counter_eq_0 : IN STD_LOGIC;
                    signal d1_OpenMAC_0_iBuf_end_xfer : IN STD_LOGIC;
                    signal d1_clock_crossing_0_s1_end_xfer : IN STD_LOGIC;
                    signal d1_cnApi_Av2Av_0_pcp_end_xfer : IN STD_LOGIC;
                    signal d1_epcs_flash_controller_0_epcs_control_port_end_xfer : IN STD_LOGIC;
                    signal d1_niosII_openMac_clock_0_in_end_xfer : IN STD_LOGIC;
                    signal d1_niosII_openMac_clock_1_in_end_xfer : IN STD_LOGIC;
                    signal d1_niosII_openMac_clock_2_in_end_xfer : IN STD_LOGIC;
                    signal d1_niosII_openMac_clock_3_in_end_xfer : IN STD_LOGIC;
                    signal d1_niosII_openMac_clock_4_in_end_xfer : IN STD_LOGIC;
                    signal d1_onchip_memory_0_s1_end_xfer : IN STD_LOGIC;
                    signal d1_pcp_cpu_jtag_debug_module_end_xfer : IN STD_LOGIC;
                    signal d1_tri_state_bridge_0_avalon_slave_end_xfer : IN STD_LOGIC;
                    signal epcs_flash_controller_0_epcs_control_port_irq_from_sa : IN STD_LOGIC;
                    signal epcs_flash_controller_0_epcs_control_port_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal incoming_tri_state_bridge_0_data : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal incoming_tri_state_bridge_0_data_with_Xs_converted_to_0 : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal jtag_uart_0_avalon_jtag_slave_irq_from_sa : IN STD_LOGIC;
                    signal niosII_openMac_clock_0_in_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal niosII_openMac_clock_0_in_waitrequest_from_sa : IN STD_LOGIC;
                    signal niosII_openMac_clock_1_in_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal niosII_openMac_clock_1_in_waitrequest_from_sa : IN STD_LOGIC;
                    signal niosII_openMac_clock_2_in_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal niosII_openMac_clock_2_in_waitrequest_from_sa : IN STD_LOGIC;
                    signal niosII_openMac_clock_3_in_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal niosII_openMac_clock_3_in_waitrequest_from_sa : IN STD_LOGIC;
                    signal niosII_openMac_clock_4_in_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal niosII_openMac_clock_4_in_waitrequest_from_sa : IN STD_LOGIC;
                    signal onchip_memory_0_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal pcp_cpu_data_master_address : IN STD_LOGIC_VECTOR (25 DOWNTO 0);
                    signal pcp_cpu_data_master_byteenable_DBC3C40_SRAM_0_avalon_tristate_slave : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal pcp_cpu_data_master_byteenable_cfi_flash_0_s1 : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal pcp_cpu_data_master_byteenable_niosII_openMac_clock_2_in : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal pcp_cpu_data_master_granted_DBC3C40_SRAM_0_avalon_tristate_slave : IN STD_LOGIC;
                    signal pcp_cpu_data_master_granted_OpenMAC_0_iBuf : IN STD_LOGIC;
                    signal pcp_cpu_data_master_granted_cfi_flash_0_s1 : IN STD_LOGIC;
                    signal pcp_cpu_data_master_granted_clock_crossing_0_s1 : IN STD_LOGIC;
                    signal pcp_cpu_data_master_granted_cnApi_Av2Av_0_pcp : IN STD_LOGIC;
                    signal pcp_cpu_data_master_granted_epcs_flash_controller_0_epcs_control_port : IN STD_LOGIC;
                    signal pcp_cpu_data_master_granted_niosII_openMac_clock_0_in : IN STD_LOGIC;
                    signal pcp_cpu_data_master_granted_niosII_openMac_clock_1_in : IN STD_LOGIC;
                    signal pcp_cpu_data_master_granted_niosII_openMac_clock_2_in : IN STD_LOGIC;
                    signal pcp_cpu_data_master_granted_niosII_openMac_clock_3_in : IN STD_LOGIC;
                    signal pcp_cpu_data_master_granted_niosII_openMac_clock_4_in : IN STD_LOGIC;
                    signal pcp_cpu_data_master_granted_onchip_memory_0_s1 : IN STD_LOGIC;
                    signal pcp_cpu_data_master_granted_pcp_cpu_jtag_debug_module : IN STD_LOGIC;
                    signal pcp_cpu_data_master_qualified_request_DBC3C40_SRAM_0_avalon_tristate_slave : IN STD_LOGIC;
                    signal pcp_cpu_data_master_qualified_request_OpenMAC_0_iBuf : IN STD_LOGIC;
                    signal pcp_cpu_data_master_qualified_request_cfi_flash_0_s1 : IN STD_LOGIC;
                    signal pcp_cpu_data_master_qualified_request_clock_crossing_0_s1 : IN STD_LOGIC;
                    signal pcp_cpu_data_master_qualified_request_cnApi_Av2Av_0_pcp : IN STD_LOGIC;
                    signal pcp_cpu_data_master_qualified_request_epcs_flash_controller_0_epcs_control_port : IN STD_LOGIC;
                    signal pcp_cpu_data_master_qualified_request_niosII_openMac_clock_0_in : IN STD_LOGIC;
                    signal pcp_cpu_data_master_qualified_request_niosII_openMac_clock_1_in : IN STD_LOGIC;
                    signal pcp_cpu_data_master_qualified_request_niosII_openMac_clock_2_in : IN STD_LOGIC;
                    signal pcp_cpu_data_master_qualified_request_niosII_openMac_clock_3_in : IN STD_LOGIC;
                    signal pcp_cpu_data_master_qualified_request_niosII_openMac_clock_4_in : IN STD_LOGIC;
                    signal pcp_cpu_data_master_qualified_request_onchip_memory_0_s1 : IN STD_LOGIC;
                    signal pcp_cpu_data_master_qualified_request_pcp_cpu_jtag_debug_module : IN STD_LOGIC;
                    signal pcp_cpu_data_master_read : IN STD_LOGIC;
                    signal pcp_cpu_data_master_read_data_valid_DBC3C40_SRAM_0_avalon_tristate_slave : IN STD_LOGIC;
                    signal pcp_cpu_data_master_read_data_valid_OpenMAC_0_iBuf : IN STD_LOGIC;
                    signal pcp_cpu_data_master_read_data_valid_cfi_flash_0_s1 : IN STD_LOGIC;
                    signal pcp_cpu_data_master_read_data_valid_clock_crossing_0_s1 : IN STD_LOGIC;
                    signal pcp_cpu_data_master_read_data_valid_clock_crossing_0_s1_shift_register : IN STD_LOGIC;
                    signal pcp_cpu_data_master_read_data_valid_cnApi_Av2Av_0_pcp : IN STD_LOGIC;
                    signal pcp_cpu_data_master_read_data_valid_epcs_flash_controller_0_epcs_control_port : IN STD_LOGIC;
                    signal pcp_cpu_data_master_read_data_valid_niosII_openMac_clock_0_in : IN STD_LOGIC;
                    signal pcp_cpu_data_master_read_data_valid_niosII_openMac_clock_1_in : IN STD_LOGIC;
                    signal pcp_cpu_data_master_read_data_valid_niosII_openMac_clock_2_in : IN STD_LOGIC;
                    signal pcp_cpu_data_master_read_data_valid_niosII_openMac_clock_3_in : IN STD_LOGIC;
                    signal pcp_cpu_data_master_read_data_valid_niosII_openMac_clock_4_in : IN STD_LOGIC;
                    signal pcp_cpu_data_master_read_data_valid_onchip_memory_0_s1 : IN STD_LOGIC;
                    signal pcp_cpu_data_master_read_data_valid_pcp_cpu_jtag_debug_module : IN STD_LOGIC;
                    signal pcp_cpu_data_master_requests_DBC3C40_SRAM_0_avalon_tristate_slave : IN STD_LOGIC;
                    signal pcp_cpu_data_master_requests_OpenMAC_0_iBuf : IN STD_LOGIC;
                    signal pcp_cpu_data_master_requests_cfi_flash_0_s1 : IN STD_LOGIC;
                    signal pcp_cpu_data_master_requests_clock_crossing_0_s1 : IN STD_LOGIC;
                    signal pcp_cpu_data_master_requests_cnApi_Av2Av_0_pcp : IN STD_LOGIC;
                    signal pcp_cpu_data_master_requests_epcs_flash_controller_0_epcs_control_port : IN STD_LOGIC;
                    signal pcp_cpu_data_master_requests_niosII_openMac_clock_0_in : IN STD_LOGIC;
                    signal pcp_cpu_data_master_requests_niosII_openMac_clock_1_in : IN STD_LOGIC;
                    signal pcp_cpu_data_master_requests_niosII_openMac_clock_2_in : IN STD_LOGIC;
                    signal pcp_cpu_data_master_requests_niosII_openMac_clock_3_in : IN STD_LOGIC;
                    signal pcp_cpu_data_master_requests_niosII_openMac_clock_4_in : IN STD_LOGIC;
                    signal pcp_cpu_data_master_requests_onchip_memory_0_s1 : IN STD_LOGIC;
                    signal pcp_cpu_data_master_requests_pcp_cpu_jtag_debug_module : IN STD_LOGIC;
                    signal pcp_cpu_data_master_write : IN STD_LOGIC;
                    signal pcp_cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal pcp_cpu_jtag_debug_module_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal registered_pcp_cpu_data_master_read_data_valid_DBC3C40_SRAM_0_avalon_tristate_slave : IN STD_LOGIC;
                    signal registered_pcp_cpu_data_master_read_data_valid_cfi_flash_0_s1 : IN STD_LOGIC;
                    signal registered_pcp_cpu_data_master_read_data_valid_onchip_memory_0_s1 : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal system_timer_s1_irq_from_sa : IN STD_LOGIC;

                 -- outputs:
                    signal pcp_cpu_data_master_address_to_slave : OUT STD_LOGIC_VECTOR (25 DOWNTO 0);
                    signal pcp_cpu_data_master_dbs_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal pcp_cpu_data_master_dbs_write_16 : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal pcp_cpu_data_master_irq : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal pcp_cpu_data_master_no_byte_enables_and_last_term : OUT STD_LOGIC;
                    signal pcp_cpu_data_master_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal pcp_cpu_data_master_waitrequest : OUT STD_LOGIC
                 );
end component pcp_cpu_data_master_arbitrator;

component pcp_cpu_instruction_master_arbitrator is 
           port (
                 -- inputs:
                    signal DBC3C40_SRAM_0_avalon_tristate_slave_wait_counter_eq_0 : IN STD_LOGIC;
                    signal cfi_flash_0_s1_wait_counter_eq_0 : IN STD_LOGIC;
                    signal cfi_flash_0_s1_wait_counter_eq_1 : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal d1_epcs_flash_controller_0_epcs_control_port_end_xfer : IN STD_LOGIC;
                    signal d1_onchip_memory_0_s1_end_xfer : IN STD_LOGIC;
                    signal d1_pcp_cpu_jtag_debug_module_end_xfer : IN STD_LOGIC;
                    signal d1_tri_state_bridge_0_avalon_slave_end_xfer : IN STD_LOGIC;
                    signal epcs_flash_controller_0_epcs_control_port_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal incoming_tri_state_bridge_0_data : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal onchip_memory_0_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal pcp_cpu_instruction_master_address : IN STD_LOGIC_VECTOR (25 DOWNTO 0);
                    signal pcp_cpu_instruction_master_granted_DBC3C40_SRAM_0_avalon_tristate_slave : IN STD_LOGIC;
                    signal pcp_cpu_instruction_master_granted_cfi_flash_0_s1 : IN STD_LOGIC;
                    signal pcp_cpu_instruction_master_granted_epcs_flash_controller_0_epcs_control_port : IN STD_LOGIC;
                    signal pcp_cpu_instruction_master_granted_onchip_memory_0_s1 : IN STD_LOGIC;
                    signal pcp_cpu_instruction_master_granted_pcp_cpu_jtag_debug_module : IN STD_LOGIC;
                    signal pcp_cpu_instruction_master_qualified_request_DBC3C40_SRAM_0_avalon_tristate_slave : IN STD_LOGIC;
                    signal pcp_cpu_instruction_master_qualified_request_cfi_flash_0_s1 : IN STD_LOGIC;
                    signal pcp_cpu_instruction_master_qualified_request_epcs_flash_controller_0_epcs_control_port : IN STD_LOGIC;
                    signal pcp_cpu_instruction_master_qualified_request_onchip_memory_0_s1 : IN STD_LOGIC;
                    signal pcp_cpu_instruction_master_qualified_request_pcp_cpu_jtag_debug_module : IN STD_LOGIC;
                    signal pcp_cpu_instruction_master_read : IN STD_LOGIC;
                    signal pcp_cpu_instruction_master_read_data_valid_DBC3C40_SRAM_0_avalon_tristate_slave : IN STD_LOGIC;
                    signal pcp_cpu_instruction_master_read_data_valid_cfi_flash_0_s1 : IN STD_LOGIC;
                    signal pcp_cpu_instruction_master_read_data_valid_epcs_flash_controller_0_epcs_control_port : IN STD_LOGIC;
                    signal pcp_cpu_instruction_master_read_data_valid_onchip_memory_0_s1 : IN STD_LOGIC;
                    signal pcp_cpu_instruction_master_read_data_valid_pcp_cpu_jtag_debug_module : IN STD_LOGIC;
                    signal pcp_cpu_instruction_master_requests_DBC3C40_SRAM_0_avalon_tristate_slave : IN STD_LOGIC;
                    signal pcp_cpu_instruction_master_requests_cfi_flash_0_s1 : IN STD_LOGIC;
                    signal pcp_cpu_instruction_master_requests_epcs_flash_controller_0_epcs_control_port : IN STD_LOGIC;
                    signal pcp_cpu_instruction_master_requests_onchip_memory_0_s1 : IN STD_LOGIC;
                    signal pcp_cpu_instruction_master_requests_pcp_cpu_jtag_debug_module : IN STD_LOGIC;
                    signal pcp_cpu_jtag_debug_module_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal pcp_cpu_instruction_master_address_to_slave : OUT STD_LOGIC_VECTOR (25 DOWNTO 0);
                    signal pcp_cpu_instruction_master_dbs_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal pcp_cpu_instruction_master_latency_counter : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal pcp_cpu_instruction_master_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal pcp_cpu_instruction_master_readdatavalid : OUT STD_LOGIC;
                    signal pcp_cpu_instruction_master_waitrequest : OUT STD_LOGIC
                 );
end component pcp_cpu_instruction_master_arbitrator;

component pcp_cpu is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal d_irq : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal d_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal d_waitrequest : IN STD_LOGIC;
                    signal i_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal i_readdatavalid : IN STD_LOGIC;
                    signal i_waitrequest : IN STD_LOGIC;
                    signal jtag_debug_module_address : IN STD_LOGIC_VECTOR (8 DOWNTO 0);
                    signal jtag_debug_module_begintransfer : IN STD_LOGIC;
                    signal jtag_debug_module_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal jtag_debug_module_debugaccess : IN STD_LOGIC;
                    signal jtag_debug_module_select : IN STD_LOGIC;
                    signal jtag_debug_module_write : IN STD_LOGIC;
                    signal jtag_debug_module_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal d_address : OUT STD_LOGIC_VECTOR (25 DOWNTO 0);
                    signal d_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal d_read : OUT STD_LOGIC;
                    signal d_write : OUT STD_LOGIC;
                    signal d_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal i_address : OUT STD_LOGIC_VECTOR (25 DOWNTO 0);
                    signal i_read : OUT STD_LOGIC;
                    signal jtag_debug_module_debugaccess_to_roms : OUT STD_LOGIC;
                    signal jtag_debug_module_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal jtag_debug_module_resetrequest : OUT STD_LOGIC
                 );
end component pcp_cpu;

component portconf_pio_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal clock_crossing_1_m1_address_to_slave : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal clock_crossing_1_m1_latency_counter : IN STD_LOGIC;
                    signal clock_crossing_1_m1_nativeaddress : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
                    signal clock_crossing_1_m1_read : IN STD_LOGIC;
                    signal clock_crossing_1_m1_write : IN STD_LOGIC;
                    signal clock_crossing_1_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal portconf_pio_s1_readdata : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal clock_crossing_1_m1_granted_portconf_pio_s1 : OUT STD_LOGIC;
                    signal clock_crossing_1_m1_qualified_request_portconf_pio_s1 : OUT STD_LOGIC;
                    signal clock_crossing_1_m1_read_data_valid_portconf_pio_s1 : OUT STD_LOGIC;
                    signal clock_crossing_1_m1_requests_portconf_pio_s1 : OUT STD_LOGIC;
                    signal d1_portconf_pio_s1_end_xfer : OUT STD_LOGIC;
                    signal portconf_pio_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal portconf_pio_s1_chipselect : OUT STD_LOGIC;
                    signal portconf_pio_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal portconf_pio_s1_reset_n : OUT STD_LOGIC;
                    signal portconf_pio_s1_write_n : OUT STD_LOGIC;
                    signal portconf_pio_s1_writedata : OUT STD_LOGIC_VECTOR (3 DOWNTO 0)
                 );
end component portconf_pio_s1_arbitrator;

component portconf_pio is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal chipselect : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal in_port : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;
                    signal write_n : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC_VECTOR (3 DOWNTO 0);

                 -- outputs:
                    signal out_port : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal readdata : OUT STD_LOGIC_VECTOR (3 DOWNTO 0)
                 );
end component portconf_pio;

component remote_update_cycloneiii_0_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal niosII_openMac_clock_4_out_address_to_slave : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal niosII_openMac_clock_4_out_nativeaddress : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
                    signal niosII_openMac_clock_4_out_read : IN STD_LOGIC;
                    signal niosII_openMac_clock_4_out_write : IN STD_LOGIC;
                    signal niosII_openMac_clock_4_out_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal remote_update_cycloneiii_0_s1_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal remote_update_cycloneiii_0_s1_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal d1_remote_update_cycloneiii_0_s1_end_xfer : OUT STD_LOGIC;
                    signal niosII_openMac_clock_4_out_granted_remote_update_cycloneiii_0_s1 : OUT STD_LOGIC;
                    signal niosII_openMac_clock_4_out_qualified_request_remote_update_cycloneiii_0_s1 : OUT STD_LOGIC;
                    signal niosII_openMac_clock_4_out_read_data_valid_remote_update_cycloneiii_0_s1 : OUT STD_LOGIC;
                    signal niosII_openMac_clock_4_out_requests_remote_update_cycloneiii_0_s1 : OUT STD_LOGIC;
                    signal remote_update_cycloneiii_0_s1_address : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
                    signal remote_update_cycloneiii_0_s1_chipselect : OUT STD_LOGIC;
                    signal remote_update_cycloneiii_0_s1_read : OUT STD_LOGIC;
                    signal remote_update_cycloneiii_0_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal remote_update_cycloneiii_0_s1_reset : OUT STD_LOGIC;
                    signal remote_update_cycloneiii_0_s1_waitrequest_from_sa : OUT STD_LOGIC;
                    signal remote_update_cycloneiii_0_s1_write : OUT STD_LOGIC;
                    signal remote_update_cycloneiii_0_s1_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
                 );
end component remote_update_cycloneiii_0_s1_arbitrator;

component remote_update_cycloneiii_0 is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
                    signal chipselect : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal waitrequest : OUT STD_LOGIC
                 );
end component remote_update_cycloneiii_0;

component sdram_0_s1_arbitrator is 
           port (
                 -- inputs:
                    signal ap_cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (25 DOWNTO 0);
                    signal ap_cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal ap_cpu_data_master_read : IN STD_LOGIC;
                    signal ap_cpu_data_master_waitrequest : IN STD_LOGIC;
                    signal ap_cpu_data_master_write : IN STD_LOGIC;
                    signal ap_cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal ap_cpu_instruction_master_address_to_slave : IN STD_LOGIC_VECTOR (25 DOWNTO 0);
                    signal ap_cpu_instruction_master_latency_counter : IN STD_LOGIC;
                    signal ap_cpu_instruction_master_read : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sdram_0_s1_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal sdram_0_s1_readdatavalid : IN STD_LOGIC;
                    signal sdram_0_s1_waitrequest : IN STD_LOGIC;

                 -- outputs:
                    signal ap_cpu_data_master_granted_sdram_0_s1 : OUT STD_LOGIC;
                    signal ap_cpu_data_master_qualified_request_sdram_0_s1 : OUT STD_LOGIC;
                    signal ap_cpu_data_master_read_data_valid_sdram_0_s1 : OUT STD_LOGIC;
                    signal ap_cpu_data_master_read_data_valid_sdram_0_s1_shift_register : OUT STD_LOGIC;
                    signal ap_cpu_data_master_requests_sdram_0_s1 : OUT STD_LOGIC;
                    signal ap_cpu_instruction_master_granted_sdram_0_s1 : OUT STD_LOGIC;
                    signal ap_cpu_instruction_master_qualified_request_sdram_0_s1 : OUT STD_LOGIC;
                    signal ap_cpu_instruction_master_read_data_valid_sdram_0_s1 : OUT STD_LOGIC;
                    signal ap_cpu_instruction_master_read_data_valid_sdram_0_s1_shift_register : OUT STD_LOGIC;
                    signal ap_cpu_instruction_master_requests_sdram_0_s1 : OUT STD_LOGIC;
                    signal d1_sdram_0_s1_end_xfer : OUT STD_LOGIC;
                    signal sdram_0_s1_address : OUT STD_LOGIC_VECTOR (21 DOWNTO 0);
                    signal sdram_0_s1_byteenable_n : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal sdram_0_s1_chipselect : OUT STD_LOGIC;
                    signal sdram_0_s1_read_n : OUT STD_LOGIC;
                    signal sdram_0_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal sdram_0_s1_reset_n : OUT STD_LOGIC;
                    signal sdram_0_s1_waitrequest_from_sa : OUT STD_LOGIC;
                    signal sdram_0_s1_write_n : OUT STD_LOGIC;
                    signal sdram_0_s1_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
                 );
end component sdram_0_s1_arbitrator;

component sdram_0 is 
           port (
                 -- inputs:
                    signal az_addr : IN STD_LOGIC_VECTOR (21 DOWNTO 0);
                    signal az_be_n : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal az_cs : IN STD_LOGIC;
                    signal az_data : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal az_rd_n : IN STD_LOGIC;
                    signal az_wr_n : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal za_data : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal za_valid : OUT STD_LOGIC;
                    signal za_waitrequest : OUT STD_LOGIC;
                    signal zs_addr : OUT STD_LOGIC_VECTOR (11 DOWNTO 0);
                    signal zs_ba : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal zs_cas_n : OUT STD_LOGIC;
                    signal zs_cke : OUT STD_LOGIC;
                    signal zs_cs_n : OUT STD_LOGIC;
                    signal zs_dq : INOUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal zs_dqm : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal zs_ras_n : OUT STD_LOGIC;
                    signal zs_we_n : OUT STD_LOGIC
                 );
end component sdram_0;

component status_led_pio_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal clock_crossing_0_m1_address_to_slave : IN STD_LOGIC_VECTOR (6 DOWNTO 0);
                    signal clock_crossing_0_m1_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal clock_crossing_0_m1_latency_counter : IN STD_LOGIC;
                    signal clock_crossing_0_m1_nativeaddress : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
                    signal clock_crossing_0_m1_read : IN STD_LOGIC;
                    signal clock_crossing_0_m1_write : IN STD_LOGIC;
                    signal clock_crossing_0_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;
                    signal status_led_pio_s1_readdata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);

                 -- outputs:
                    signal clock_crossing_0_m1_granted_status_led_pio_s1 : OUT STD_LOGIC;
                    signal clock_crossing_0_m1_qualified_request_status_led_pio_s1 : OUT STD_LOGIC;
                    signal clock_crossing_0_m1_read_data_valid_status_led_pio_s1 : OUT STD_LOGIC;
                    signal clock_crossing_0_m1_requests_status_led_pio_s1 : OUT STD_LOGIC;
                    signal d1_status_led_pio_s1_end_xfer : OUT STD_LOGIC;
                    signal status_led_pio_s1_address : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal status_led_pio_s1_chipselect : OUT STD_LOGIC;
                    signal status_led_pio_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal status_led_pio_s1_reset_n : OUT STD_LOGIC;
                    signal status_led_pio_s1_write_n : OUT STD_LOGIC;
                    signal status_led_pio_s1_writedata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
                 );
end component status_led_pio_s1_arbitrator;

component status_led_pio is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal chipselect : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal write_n : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);

                 -- outputs:
                    signal out_port : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal readdata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
                 );
end component status_led_pio;

component sync_irq_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal clock_crossing_1_m1_address_to_slave : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal clock_crossing_1_m1_latency_counter : IN STD_LOGIC;
                    signal clock_crossing_1_m1_nativeaddress : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
                    signal clock_crossing_1_m1_read : IN STD_LOGIC;
                    signal clock_crossing_1_m1_write : IN STD_LOGIC;
                    signal clock_crossing_1_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;
                    signal sync_irq_s1_irq : IN STD_LOGIC;
                    signal sync_irq_s1_readdata : IN STD_LOGIC;

                 -- outputs:
                    signal clock_crossing_1_m1_granted_sync_irq_s1 : OUT STD_LOGIC;
                    signal clock_crossing_1_m1_qualified_request_sync_irq_s1 : OUT STD_LOGIC;
                    signal clock_crossing_1_m1_read_data_valid_sync_irq_s1 : OUT STD_LOGIC;
                    signal clock_crossing_1_m1_requests_sync_irq_s1 : OUT STD_LOGIC;
                    signal d1_sync_irq_s1_end_xfer : OUT STD_LOGIC;
                    signal sync_irq_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal sync_irq_s1_chipselect : OUT STD_LOGIC;
                    signal sync_irq_s1_irq_from_sa : OUT STD_LOGIC;
                    signal sync_irq_s1_readdata_from_sa : OUT STD_LOGIC;
                    signal sync_irq_s1_reset_n : OUT STD_LOGIC;
                    signal sync_irq_s1_write_n : OUT STD_LOGIC;
                    signal sync_irq_s1_writedata : OUT STD_LOGIC
                 );
end component sync_irq_s1_arbitrator;

component sync_irq is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal chipselect : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal in_port : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal write_n : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC;

                 -- outputs:
                    signal irq : OUT STD_LOGIC;
                    signal readdata : OUT STD_LOGIC
                 );
end component sync_irq;

component sysid_control_slave_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal clock_crossing_0_m1_address_to_slave : IN STD_LOGIC_VECTOR (6 DOWNTO 0);
                    signal clock_crossing_0_m1_latency_counter : IN STD_LOGIC;
                    signal clock_crossing_0_m1_nativeaddress : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
                    signal clock_crossing_0_m1_read : IN STD_LOGIC;
                    signal clock_crossing_0_m1_write : IN STD_LOGIC;
                    signal clock_crossing_1_m1_address_to_slave : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal clock_crossing_1_m1_latency_counter : IN STD_LOGIC;
                    signal clock_crossing_1_m1_nativeaddress : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
                    signal clock_crossing_1_m1_read : IN STD_LOGIC;
                    signal clock_crossing_1_m1_write : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sysid_control_slave_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal clock_crossing_0_m1_granted_sysid_control_slave : OUT STD_LOGIC;
                    signal clock_crossing_0_m1_qualified_request_sysid_control_slave : OUT STD_LOGIC;
                    signal clock_crossing_0_m1_read_data_valid_sysid_control_slave : OUT STD_LOGIC;
                    signal clock_crossing_0_m1_requests_sysid_control_slave : OUT STD_LOGIC;
                    signal clock_crossing_1_m1_granted_sysid_control_slave : OUT STD_LOGIC;
                    signal clock_crossing_1_m1_qualified_request_sysid_control_slave : OUT STD_LOGIC;
                    signal clock_crossing_1_m1_read_data_valid_sysid_control_slave : OUT STD_LOGIC;
                    signal clock_crossing_1_m1_requests_sysid_control_slave : OUT STD_LOGIC;
                    signal d1_sysid_control_slave_end_xfer : OUT STD_LOGIC;
                    signal sysid_control_slave_address : OUT STD_LOGIC;
                    signal sysid_control_slave_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
                 );
end component sysid_control_slave_arbitrator;

component sysid is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC;

                 -- outputs:
                    signal readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
                 );
end component sysid;

component system_timer_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal clock_crossing_0_m1_address_to_slave : IN STD_LOGIC_VECTOR (6 DOWNTO 0);
                    signal clock_crossing_0_m1_latency_counter : IN STD_LOGIC;
                    signal clock_crossing_0_m1_nativeaddress : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
                    signal clock_crossing_0_m1_read : IN STD_LOGIC;
                    signal clock_crossing_0_m1_write : IN STD_LOGIC;
                    signal clock_crossing_0_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;
                    signal system_timer_s1_irq : IN STD_LOGIC;
                    signal system_timer_s1_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

                 -- outputs:
                    signal clock_crossing_0_m1_granted_system_timer_s1 : OUT STD_LOGIC;
                    signal clock_crossing_0_m1_qualified_request_system_timer_s1 : OUT STD_LOGIC;
                    signal clock_crossing_0_m1_read_data_valid_system_timer_s1 : OUT STD_LOGIC;
                    signal clock_crossing_0_m1_requests_system_timer_s1 : OUT STD_LOGIC;
                    signal d1_system_timer_s1_end_xfer : OUT STD_LOGIC;
                    signal system_timer_s1_address : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal system_timer_s1_chipselect : OUT STD_LOGIC;
                    signal system_timer_s1_irq_from_sa : OUT STD_LOGIC;
                    signal system_timer_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal system_timer_s1_reset_n : OUT STD_LOGIC;
                    signal system_timer_s1_write_n : OUT STD_LOGIC;
                    signal system_timer_s1_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
                 );
end component system_timer_s1_arbitrator;

component system_timer is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal chipselect : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal write_n : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

                 -- outputs:
                    signal irq : OUT STD_LOGIC;
                    signal readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
                 );
end component system_timer;

component system_timer_ap_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal clock_crossing_1_m1_address_to_slave : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal clock_crossing_1_m1_latency_counter : IN STD_LOGIC;
                    signal clock_crossing_1_m1_nativeaddress : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
                    signal clock_crossing_1_m1_read : IN STD_LOGIC;
                    signal clock_crossing_1_m1_write : IN STD_LOGIC;
                    signal clock_crossing_1_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;
                    signal system_timer_ap_s1_irq : IN STD_LOGIC;
                    signal system_timer_ap_s1_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

                 -- outputs:
                    signal clock_crossing_1_m1_granted_system_timer_ap_s1 : OUT STD_LOGIC;
                    signal clock_crossing_1_m1_qualified_request_system_timer_ap_s1 : OUT STD_LOGIC;
                    signal clock_crossing_1_m1_read_data_valid_system_timer_ap_s1 : OUT STD_LOGIC;
                    signal clock_crossing_1_m1_requests_system_timer_ap_s1 : OUT STD_LOGIC;
                    signal d1_system_timer_ap_s1_end_xfer : OUT STD_LOGIC;
                    signal system_timer_ap_s1_address : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal system_timer_ap_s1_chipselect : OUT STD_LOGIC;
                    signal system_timer_ap_s1_irq_from_sa : OUT STD_LOGIC;
                    signal system_timer_ap_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal system_timer_ap_s1_reset_n : OUT STD_LOGIC;
                    signal system_timer_ap_s1_write_n : OUT STD_LOGIC;
                    signal system_timer_ap_s1_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
                 );
end component system_timer_ap_s1_arbitrator;

component system_timer_ap is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal chipselect : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal write_n : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

                 -- outputs:
                    signal irq : OUT STD_LOGIC;
                    signal readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
                 );
end component system_timer_ap;

component tri_state_bridge_0_avalon_slave_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal pcp_cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (25 DOWNTO 0);
                    signal pcp_cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal pcp_cpu_data_master_dbs_address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal pcp_cpu_data_master_dbs_write_16 : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal pcp_cpu_data_master_no_byte_enables_and_last_term : IN STD_LOGIC;
                    signal pcp_cpu_data_master_read : IN STD_LOGIC;
                    signal pcp_cpu_data_master_write : IN STD_LOGIC;
                    signal pcp_cpu_instruction_master_address_to_slave : IN STD_LOGIC_VECTOR (25 DOWNTO 0);
                    signal pcp_cpu_instruction_master_dbs_address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal pcp_cpu_instruction_master_latency_counter : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal pcp_cpu_instruction_master_read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal DBC3C40_SRAM_0_avalon_tristate_slave_wait_counter_eq_0 : OUT STD_LOGIC;
                    signal ben_to_the_DBC3C40_SRAM_0 : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal cfi_flash_0_s1_wait_counter_eq_0 : OUT STD_LOGIC;
                    signal cfi_flash_0_s1_wait_counter_eq_1 : OUT STD_LOGIC;
                    signal d1_tri_state_bridge_0_avalon_slave_end_xfer : OUT STD_LOGIC;
                    signal incoming_tri_state_bridge_0_data : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal incoming_tri_state_bridge_0_data_with_Xs_converted_to_0 : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal ncs_to_the_DBC3C40_SRAM_0 : OUT STD_LOGIC;
                    signal pcp_cpu_data_master_byteenable_DBC3C40_SRAM_0_avalon_tristate_slave : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal pcp_cpu_data_master_byteenable_cfi_flash_0_s1 : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal pcp_cpu_data_master_granted_DBC3C40_SRAM_0_avalon_tristate_slave : OUT STD_LOGIC;
                    signal pcp_cpu_data_master_granted_cfi_flash_0_s1 : OUT STD_LOGIC;
                    signal pcp_cpu_data_master_qualified_request_DBC3C40_SRAM_0_avalon_tristate_slave : OUT STD_LOGIC;
                    signal pcp_cpu_data_master_qualified_request_cfi_flash_0_s1 : OUT STD_LOGIC;
                    signal pcp_cpu_data_master_read_data_valid_DBC3C40_SRAM_0_avalon_tristate_slave : OUT STD_LOGIC;
                    signal pcp_cpu_data_master_read_data_valid_cfi_flash_0_s1 : OUT STD_LOGIC;
                    signal pcp_cpu_data_master_requests_DBC3C40_SRAM_0_avalon_tristate_slave : OUT STD_LOGIC;
                    signal pcp_cpu_data_master_requests_cfi_flash_0_s1 : OUT STD_LOGIC;
                    signal pcp_cpu_instruction_master_granted_DBC3C40_SRAM_0_avalon_tristate_slave : OUT STD_LOGIC;
                    signal pcp_cpu_instruction_master_granted_cfi_flash_0_s1 : OUT STD_LOGIC;
                    signal pcp_cpu_instruction_master_qualified_request_DBC3C40_SRAM_0_avalon_tristate_slave : OUT STD_LOGIC;
                    signal pcp_cpu_instruction_master_qualified_request_cfi_flash_0_s1 : OUT STD_LOGIC;
                    signal pcp_cpu_instruction_master_read_data_valid_DBC3C40_SRAM_0_avalon_tristate_slave : OUT STD_LOGIC;
                    signal pcp_cpu_instruction_master_read_data_valid_cfi_flash_0_s1 : OUT STD_LOGIC;
                    signal pcp_cpu_instruction_master_requests_DBC3C40_SRAM_0_avalon_tristate_slave : OUT STD_LOGIC;
                    signal pcp_cpu_instruction_master_requests_cfi_flash_0_s1 : OUT STD_LOGIC;
                    signal registered_pcp_cpu_data_master_read_data_valid_DBC3C40_SRAM_0_avalon_tristate_slave : OUT STD_LOGIC;
                    signal registered_pcp_cpu_data_master_read_data_valid_cfi_flash_0_s1 : OUT STD_LOGIC;
                    signal select_n_to_the_cfi_flash_0 : OUT STD_LOGIC;
                    signal tri_state_bridge_0_address : OUT STD_LOGIC_VECTOR (22 DOWNTO 0);
                    signal tri_state_bridge_0_data : INOUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal tri_state_bridge_0_readn : OUT STD_LOGIC;
                    signal tri_state_bridge_0_writen : OUT STD_LOGIC
                 );
end component tri_state_bridge_0_avalon_slave_arbitrator;

component tri_state_bridge_0 is 
end component tri_state_bridge_0;

component tri_state_bridge_0_bridge_arbitrator is 
end component tri_state_bridge_0_bridge_arbitrator;

component niosII_openMac_reset_clk50Meg_domain_synch_module is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC
                 );
end component niosII_openMac_reset_clk50Meg_domain_synch_module;

component niosII_openMac_reset_clk90Meg_domain_synch_module is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC
                 );
end component niosII_openMac_reset_clk90Meg_domain_synch_module;

component niosII_openMac_reset_clk_0_domain_synch_module is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC
                 );
end component niosII_openMac_reset_clk_0_domain_synch_module;

component niosII_openMac_reset_clk25Meg_domain_synch_module is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC
                 );
end component niosII_openMac_reset_clk25Meg_domain_synch_module;

                signal DBC3C40_SRAM_0_avalon_tristate_slave_wait_counter_eq_0 :  STD_LOGIC;
                signal OpenMAC_0_CMP_address :  STD_LOGIC;
                signal OpenMAC_0_CMP_byteenable_n :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal OpenMAC_0_CMP_chipselect :  STD_LOGIC;
                signal OpenMAC_0_CMP_irq :  STD_LOGIC;
                signal OpenMAC_0_CMP_irq_from_sa :  STD_LOGIC;
                signal OpenMAC_0_CMP_read_n :  STD_LOGIC;
                signal OpenMAC_0_CMP_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal OpenMAC_0_CMP_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal OpenMAC_0_CMP_reset_n :  STD_LOGIC;
                signal OpenMAC_0_CMP_write_n :  STD_LOGIC;
                signal OpenMAC_0_CMP_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal OpenMAC_0_REG_address :  STD_LOGIC_VECTOR (11 DOWNTO 0);
                signal OpenMAC_0_REG_byteenable_n :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal OpenMAC_0_REG_chipselect :  STD_LOGIC;
                signal OpenMAC_0_REG_irq :  STD_LOGIC;
                signal OpenMAC_0_REG_irq_from_sa :  STD_LOGIC;
                signal OpenMAC_0_REG_read_n :  STD_LOGIC;
                signal OpenMAC_0_REG_readdata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal OpenMAC_0_REG_readdata_from_sa :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal OpenMAC_0_REG_write_n :  STD_LOGIC;
                signal OpenMAC_0_REG_writedata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal OpenMAC_0_iBuf_address :  STD_LOGIC_VECTOR (12 DOWNTO 0);
                signal OpenMAC_0_iBuf_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal OpenMAC_0_iBuf_chipselect :  STD_LOGIC;
                signal OpenMAC_0_iBuf_read_n :  STD_LOGIC;
                signal OpenMAC_0_iBuf_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal OpenMAC_0_iBuf_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal OpenMAC_0_iBuf_wait_counter_eq_0 :  STD_LOGIC;
                signal OpenMAC_0_iBuf_write_n :  STD_LOGIC;
                signal OpenMAC_0_iBuf_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal altpll_0_pll_slave_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal altpll_0_pll_slave_read :  STD_LOGIC;
                signal altpll_0_pll_slave_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal altpll_0_pll_slave_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal altpll_0_pll_slave_reset :  STD_LOGIC;
                signal altpll_0_pll_slave_write :  STD_LOGIC;
                signal altpll_0_pll_slave_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal ap_cpu_data_master_address :  STD_LOGIC_VECTOR (25 DOWNTO 0);
                signal ap_cpu_data_master_address_to_slave :  STD_LOGIC_VECTOR (25 DOWNTO 0);
                signal ap_cpu_data_master_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal ap_cpu_data_master_debugaccess :  STD_LOGIC;
                signal ap_cpu_data_master_granted_ap_cpu_jtag_debug_module :  STD_LOGIC;
                signal ap_cpu_data_master_granted_clock_crossing_1_s1 :  STD_LOGIC;
                signal ap_cpu_data_master_granted_cnApi_Av2Av_0_ap :  STD_LOGIC;
                signal ap_cpu_data_master_granted_jtag_uart_1_avalon_jtag_slave :  STD_LOGIC;
                signal ap_cpu_data_master_granted_sdram_0_s1 :  STD_LOGIC;
                signal ap_cpu_data_master_irq :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal ap_cpu_data_master_qualified_request_ap_cpu_jtag_debug_module :  STD_LOGIC;
                signal ap_cpu_data_master_qualified_request_clock_crossing_1_s1 :  STD_LOGIC;
                signal ap_cpu_data_master_qualified_request_cnApi_Av2Av_0_ap :  STD_LOGIC;
                signal ap_cpu_data_master_qualified_request_jtag_uart_1_avalon_jtag_slave :  STD_LOGIC;
                signal ap_cpu_data_master_qualified_request_sdram_0_s1 :  STD_LOGIC;
                signal ap_cpu_data_master_read :  STD_LOGIC;
                signal ap_cpu_data_master_read_data_valid_ap_cpu_jtag_debug_module :  STD_LOGIC;
                signal ap_cpu_data_master_read_data_valid_clock_crossing_1_s1 :  STD_LOGIC;
                signal ap_cpu_data_master_read_data_valid_clock_crossing_1_s1_shift_register :  STD_LOGIC;
                signal ap_cpu_data_master_read_data_valid_cnApi_Av2Av_0_ap :  STD_LOGIC;
                signal ap_cpu_data_master_read_data_valid_jtag_uart_1_avalon_jtag_slave :  STD_LOGIC;
                signal ap_cpu_data_master_read_data_valid_sdram_0_s1 :  STD_LOGIC;
                signal ap_cpu_data_master_read_data_valid_sdram_0_s1_shift_register :  STD_LOGIC;
                signal ap_cpu_data_master_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal ap_cpu_data_master_requests_ap_cpu_jtag_debug_module :  STD_LOGIC;
                signal ap_cpu_data_master_requests_clock_crossing_1_s1 :  STD_LOGIC;
                signal ap_cpu_data_master_requests_cnApi_Av2Av_0_ap :  STD_LOGIC;
                signal ap_cpu_data_master_requests_jtag_uart_1_avalon_jtag_slave :  STD_LOGIC;
                signal ap_cpu_data_master_requests_sdram_0_s1 :  STD_LOGIC;
                signal ap_cpu_data_master_waitrequest :  STD_LOGIC;
                signal ap_cpu_data_master_write :  STD_LOGIC;
                signal ap_cpu_data_master_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal ap_cpu_instruction_master_address :  STD_LOGIC_VECTOR (25 DOWNTO 0);
                signal ap_cpu_instruction_master_address_to_slave :  STD_LOGIC_VECTOR (25 DOWNTO 0);
                signal ap_cpu_instruction_master_granted_ap_cpu_jtag_debug_module :  STD_LOGIC;
                signal ap_cpu_instruction_master_granted_sdram_0_s1 :  STD_LOGIC;
                signal ap_cpu_instruction_master_latency_counter :  STD_LOGIC;
                signal ap_cpu_instruction_master_qualified_request_ap_cpu_jtag_debug_module :  STD_LOGIC;
                signal ap_cpu_instruction_master_qualified_request_sdram_0_s1 :  STD_LOGIC;
                signal ap_cpu_instruction_master_read :  STD_LOGIC;
                signal ap_cpu_instruction_master_read_data_valid_ap_cpu_jtag_debug_module :  STD_LOGIC;
                signal ap_cpu_instruction_master_read_data_valid_sdram_0_s1 :  STD_LOGIC;
                signal ap_cpu_instruction_master_read_data_valid_sdram_0_s1_shift_register :  STD_LOGIC;
                signal ap_cpu_instruction_master_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal ap_cpu_instruction_master_readdatavalid :  STD_LOGIC;
                signal ap_cpu_instruction_master_requests_ap_cpu_jtag_debug_module :  STD_LOGIC;
                signal ap_cpu_instruction_master_requests_sdram_0_s1 :  STD_LOGIC;
                signal ap_cpu_instruction_master_waitrequest :  STD_LOGIC;
                signal ap_cpu_jtag_debug_module_address :  STD_LOGIC_VECTOR (8 DOWNTO 0);
                signal ap_cpu_jtag_debug_module_begintransfer :  STD_LOGIC;
                signal ap_cpu_jtag_debug_module_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal ap_cpu_jtag_debug_module_chipselect :  STD_LOGIC;
                signal ap_cpu_jtag_debug_module_debugaccess :  STD_LOGIC;
                signal ap_cpu_jtag_debug_module_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal ap_cpu_jtag_debug_module_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal ap_cpu_jtag_debug_module_reset_n :  STD_LOGIC;
                signal ap_cpu_jtag_debug_module_resetrequest :  STD_LOGIC;
                signal ap_cpu_jtag_debug_module_resetrequest_from_sa :  STD_LOGIC;
                signal ap_cpu_jtag_debug_module_write :  STD_LOGIC;
                signal ap_cpu_jtag_debug_module_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal button_pio_s1_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal button_pio_s1_readdata :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal button_pio_s1_readdata_from_sa :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal button_pio_s1_reset_n :  STD_LOGIC;
                signal cfi_flash_0_s1_wait_counter_eq_0 :  STD_LOGIC;
                signal cfi_flash_0_s1_wait_counter_eq_1 :  STD_LOGIC;
                signal clk25Meg_reset_n :  STD_LOGIC;
                signal clk50Meg_reset_n :  STD_LOGIC;
                signal clk90Meg_reset_n :  STD_LOGIC;
                signal clk_0_reset_n :  STD_LOGIC;
                signal clock_crossing_0_m1_address :  STD_LOGIC_VECTOR (6 DOWNTO 0);
                signal clock_crossing_0_m1_address_to_slave :  STD_LOGIC_VECTOR (6 DOWNTO 0);
                signal clock_crossing_0_m1_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal clock_crossing_0_m1_endofpacket :  STD_LOGIC;
                signal clock_crossing_0_m1_granted_button_pio_s1 :  STD_LOGIC;
                signal clock_crossing_0_m1_granted_irq_gen_s1 :  STD_LOGIC;
                signal clock_crossing_0_m1_granted_status_led_pio_s1 :  STD_LOGIC;
                signal clock_crossing_0_m1_granted_sysid_control_slave :  STD_LOGIC;
                signal clock_crossing_0_m1_granted_system_timer_s1 :  STD_LOGIC;
                signal clock_crossing_0_m1_latency_counter :  STD_LOGIC;
                signal clock_crossing_0_m1_nativeaddress :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal clock_crossing_0_m1_qualified_request_button_pio_s1 :  STD_LOGIC;
                signal clock_crossing_0_m1_qualified_request_irq_gen_s1 :  STD_LOGIC;
                signal clock_crossing_0_m1_qualified_request_status_led_pio_s1 :  STD_LOGIC;
                signal clock_crossing_0_m1_qualified_request_sysid_control_slave :  STD_LOGIC;
                signal clock_crossing_0_m1_qualified_request_system_timer_s1 :  STD_LOGIC;
                signal clock_crossing_0_m1_read :  STD_LOGIC;
                signal clock_crossing_0_m1_read_data_valid_button_pio_s1 :  STD_LOGIC;
                signal clock_crossing_0_m1_read_data_valid_irq_gen_s1 :  STD_LOGIC;
                signal clock_crossing_0_m1_read_data_valid_status_led_pio_s1 :  STD_LOGIC;
                signal clock_crossing_0_m1_read_data_valid_sysid_control_slave :  STD_LOGIC;
                signal clock_crossing_0_m1_read_data_valid_system_timer_s1 :  STD_LOGIC;
                signal clock_crossing_0_m1_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal clock_crossing_0_m1_readdatavalid :  STD_LOGIC;
                signal clock_crossing_0_m1_requests_button_pio_s1 :  STD_LOGIC;
                signal clock_crossing_0_m1_requests_irq_gen_s1 :  STD_LOGIC;
                signal clock_crossing_0_m1_requests_status_led_pio_s1 :  STD_LOGIC;
                signal clock_crossing_0_m1_requests_sysid_control_slave :  STD_LOGIC;
                signal clock_crossing_0_m1_requests_system_timer_s1 :  STD_LOGIC;
                signal clock_crossing_0_m1_reset_n :  STD_LOGIC;
                signal clock_crossing_0_m1_waitrequest :  STD_LOGIC;
                signal clock_crossing_0_m1_write :  STD_LOGIC;
                signal clock_crossing_0_m1_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal clock_crossing_0_s1_address :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal clock_crossing_0_s1_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal clock_crossing_0_s1_endofpacket :  STD_LOGIC;
                signal clock_crossing_0_s1_endofpacket_from_sa :  STD_LOGIC;
                signal clock_crossing_0_s1_nativeaddress :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal clock_crossing_0_s1_read :  STD_LOGIC;
                signal clock_crossing_0_s1_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal clock_crossing_0_s1_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal clock_crossing_0_s1_readdatavalid :  STD_LOGIC;
                signal clock_crossing_0_s1_reset_n :  STD_LOGIC;
                signal clock_crossing_0_s1_waitrequest :  STD_LOGIC;
                signal clock_crossing_0_s1_waitrequest_from_sa :  STD_LOGIC;
                signal clock_crossing_0_s1_write :  STD_LOGIC;
                signal clock_crossing_0_s1_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal clock_crossing_1_m1_address :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal clock_crossing_1_m1_address_to_slave :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal clock_crossing_1_m1_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal clock_crossing_1_m1_endofpacket :  STD_LOGIC;
                signal clock_crossing_1_m1_granted_digio_pio_s1 :  STD_LOGIC;
                signal clock_crossing_1_m1_granted_node_switch_pio_s1 :  STD_LOGIC;
                signal clock_crossing_1_m1_granted_portconf_pio_s1 :  STD_LOGIC;
                signal clock_crossing_1_m1_granted_sync_irq_s1 :  STD_LOGIC;
                signal clock_crossing_1_m1_granted_sysid_control_slave :  STD_LOGIC;
                signal clock_crossing_1_m1_granted_system_timer_ap_s1 :  STD_LOGIC;
                signal clock_crossing_1_m1_latency_counter :  STD_LOGIC;
                signal clock_crossing_1_m1_nativeaddress :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal clock_crossing_1_m1_qualified_request_digio_pio_s1 :  STD_LOGIC;
                signal clock_crossing_1_m1_qualified_request_node_switch_pio_s1 :  STD_LOGIC;
                signal clock_crossing_1_m1_qualified_request_portconf_pio_s1 :  STD_LOGIC;
                signal clock_crossing_1_m1_qualified_request_sync_irq_s1 :  STD_LOGIC;
                signal clock_crossing_1_m1_qualified_request_sysid_control_slave :  STD_LOGIC;
                signal clock_crossing_1_m1_qualified_request_system_timer_ap_s1 :  STD_LOGIC;
                signal clock_crossing_1_m1_read :  STD_LOGIC;
                signal clock_crossing_1_m1_read_data_valid_digio_pio_s1 :  STD_LOGIC;
                signal clock_crossing_1_m1_read_data_valid_node_switch_pio_s1 :  STD_LOGIC;
                signal clock_crossing_1_m1_read_data_valid_portconf_pio_s1 :  STD_LOGIC;
                signal clock_crossing_1_m1_read_data_valid_sync_irq_s1 :  STD_LOGIC;
                signal clock_crossing_1_m1_read_data_valid_sysid_control_slave :  STD_LOGIC;
                signal clock_crossing_1_m1_read_data_valid_system_timer_ap_s1 :  STD_LOGIC;
                signal clock_crossing_1_m1_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal clock_crossing_1_m1_readdatavalid :  STD_LOGIC;
                signal clock_crossing_1_m1_requests_digio_pio_s1 :  STD_LOGIC;
                signal clock_crossing_1_m1_requests_node_switch_pio_s1 :  STD_LOGIC;
                signal clock_crossing_1_m1_requests_portconf_pio_s1 :  STD_LOGIC;
                signal clock_crossing_1_m1_requests_sync_irq_s1 :  STD_LOGIC;
                signal clock_crossing_1_m1_requests_sysid_control_slave :  STD_LOGIC;
                signal clock_crossing_1_m1_requests_system_timer_ap_s1 :  STD_LOGIC;
                signal clock_crossing_1_m1_reset_n :  STD_LOGIC;
                signal clock_crossing_1_m1_waitrequest :  STD_LOGIC;
                signal clock_crossing_1_m1_write :  STD_LOGIC;
                signal clock_crossing_1_m1_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal clock_crossing_1_s1_address :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal clock_crossing_1_s1_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal clock_crossing_1_s1_endofpacket :  STD_LOGIC;
                signal clock_crossing_1_s1_endofpacket_from_sa :  STD_LOGIC;
                signal clock_crossing_1_s1_nativeaddress :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal clock_crossing_1_s1_read :  STD_LOGIC;
                signal clock_crossing_1_s1_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal clock_crossing_1_s1_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal clock_crossing_1_s1_readdatavalid :  STD_LOGIC;
                signal clock_crossing_1_s1_reset_n :  STD_LOGIC;
                signal clock_crossing_1_s1_waitrequest :  STD_LOGIC;
                signal clock_crossing_1_s1_waitrequest_from_sa :  STD_LOGIC;
                signal clock_crossing_1_s1_write :  STD_LOGIC;
                signal clock_crossing_1_s1_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal cnApi_Av2Av_0_ap_address :  STD_LOGIC_VECTOR (14 DOWNTO 0);
                signal cnApi_Av2Av_0_ap_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal cnApi_Av2Av_0_ap_chipselect :  STD_LOGIC;
                signal cnApi_Av2Av_0_ap_read :  STD_LOGIC;
                signal cnApi_Av2Av_0_ap_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal cnApi_Av2Av_0_ap_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal cnApi_Av2Av_0_ap_reset :  STD_LOGIC;
                signal cnApi_Av2Av_0_ap_wait_counter_eq_0 :  STD_LOGIC;
                signal cnApi_Av2Av_0_ap_write :  STD_LOGIC;
                signal cnApi_Av2Av_0_ap_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal cnApi_Av2Av_0_pcp_address :  STD_LOGIC_VECTOR (14 DOWNTO 0);
                signal cnApi_Av2Av_0_pcp_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal cnApi_Av2Av_0_pcp_chipselect :  STD_LOGIC;
                signal cnApi_Av2Av_0_pcp_read :  STD_LOGIC;
                signal cnApi_Av2Av_0_pcp_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal cnApi_Av2Av_0_pcp_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal cnApi_Av2Av_0_pcp_reset :  STD_LOGIC;
                signal cnApi_Av2Av_0_pcp_wait_counter_eq_0 :  STD_LOGIC;
                signal cnApi_Av2Av_0_pcp_write :  STD_LOGIC;
                signal cnApi_Av2Av_0_pcp_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal d1_OpenMAC_0_CMP_end_xfer :  STD_LOGIC;
                signal d1_OpenMAC_0_REG_end_xfer :  STD_LOGIC;
                signal d1_OpenMAC_0_iBuf_end_xfer :  STD_LOGIC;
                signal d1_altpll_0_pll_slave_end_xfer :  STD_LOGIC;
                signal d1_ap_cpu_jtag_debug_module_end_xfer :  STD_LOGIC;
                signal d1_button_pio_s1_end_xfer :  STD_LOGIC;
                signal d1_clock_crossing_0_s1_end_xfer :  STD_LOGIC;
                signal d1_clock_crossing_1_s1_end_xfer :  STD_LOGIC;
                signal d1_cnApi_Av2Av_0_ap_end_xfer :  STD_LOGIC;
                signal d1_cnApi_Av2Av_0_pcp_end_xfer :  STD_LOGIC;
                signal d1_digio_pio_s1_end_xfer :  STD_LOGIC;
                signal d1_epcs_flash_controller_0_epcs_control_port_end_xfer :  STD_LOGIC;
                signal d1_irq_gen_s1_end_xfer :  STD_LOGIC;
                signal d1_jtag_uart_0_avalon_jtag_slave_end_xfer :  STD_LOGIC;
                signal d1_jtag_uart_1_avalon_jtag_slave_end_xfer :  STD_LOGIC;
                signal d1_niosII_openMac_clock_0_in_end_xfer :  STD_LOGIC;
                signal d1_niosII_openMac_clock_1_in_end_xfer :  STD_LOGIC;
                signal d1_niosII_openMac_clock_2_in_end_xfer :  STD_LOGIC;
                signal d1_niosII_openMac_clock_3_in_end_xfer :  STD_LOGIC;
                signal d1_niosII_openMac_clock_4_in_end_xfer :  STD_LOGIC;
                signal d1_node_switch_pio_s1_end_xfer :  STD_LOGIC;
                signal d1_onchip_memory_0_s1_end_xfer :  STD_LOGIC;
                signal d1_pcp_cpu_jtag_debug_module_end_xfer :  STD_LOGIC;
                signal d1_portconf_pio_s1_end_xfer :  STD_LOGIC;
                signal d1_remote_update_cycloneiii_0_s1_end_xfer :  STD_LOGIC;
                signal d1_sdram_0_s1_end_xfer :  STD_LOGIC;
                signal d1_status_led_pio_s1_end_xfer :  STD_LOGIC;
                signal d1_sync_irq_s1_end_xfer :  STD_LOGIC;
                signal d1_sysid_control_slave_end_xfer :  STD_LOGIC;
                signal d1_system_timer_ap_s1_end_xfer :  STD_LOGIC;
                signal d1_system_timer_s1_end_xfer :  STD_LOGIC;
                signal d1_tri_state_bridge_0_avalon_slave_end_xfer :  STD_LOGIC;
                signal digio_pio_s1_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal digio_pio_s1_chipselect :  STD_LOGIC;
                signal digio_pio_s1_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal digio_pio_s1_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal digio_pio_s1_reset_n :  STD_LOGIC;
                signal digio_pio_s1_write_n :  STD_LOGIC;
                signal digio_pio_s1_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal epcs_flash_controller_0_epcs_control_port_address :  STD_LOGIC_VECTOR (8 DOWNTO 0);
                signal epcs_flash_controller_0_epcs_control_port_chipselect :  STD_LOGIC;
                signal epcs_flash_controller_0_epcs_control_port_dataavailable :  STD_LOGIC;
                signal epcs_flash_controller_0_epcs_control_port_dataavailable_from_sa :  STD_LOGIC;
                signal epcs_flash_controller_0_epcs_control_port_endofpacket :  STD_LOGIC;
                signal epcs_flash_controller_0_epcs_control_port_endofpacket_from_sa :  STD_LOGIC;
                signal epcs_flash_controller_0_epcs_control_port_irq :  STD_LOGIC;
                signal epcs_flash_controller_0_epcs_control_port_irq_from_sa :  STD_LOGIC;
                signal epcs_flash_controller_0_epcs_control_port_read_n :  STD_LOGIC;
                signal epcs_flash_controller_0_epcs_control_port_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal epcs_flash_controller_0_epcs_control_port_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal epcs_flash_controller_0_epcs_control_port_readyfordata :  STD_LOGIC;
                signal epcs_flash_controller_0_epcs_control_port_readyfordata_from_sa :  STD_LOGIC;
                signal epcs_flash_controller_0_epcs_control_port_reset_n :  STD_LOGIC;
                signal epcs_flash_controller_0_epcs_control_port_write_n :  STD_LOGIC;
                signal epcs_flash_controller_0_epcs_control_port_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal incoming_tri_state_bridge_0_data :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal incoming_tri_state_bridge_0_data_with_Xs_converted_to_0 :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal internal_ben_to_the_DBC3C40_SRAM_0 :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal internal_clk25Meg :  STD_LOGIC;
                signal internal_clk50Meg :  STD_LOGIC;
                signal internal_clk90Meg :  STD_LOGIC;
                signal internal_dclk_from_the_epcs_flash_controller_0 :  STD_LOGIC;
                signal internal_locked_from_the_altpll_0 :  STD_LOGIC;
                signal internal_mii_Clk_from_the_OpenMAC_0 :  STD_LOGIC;
                signal internal_mii_Do_from_the_OpenMAC_0 :  STD_LOGIC;
                signal internal_mii_Doe_from_the_OpenMAC_0 :  STD_LOGIC;
                signal internal_mii_nResetOut_from_the_OpenMAC_0 :  STD_LOGIC;
                signal internal_ncs_to_the_DBC3C40_SRAM_0 :  STD_LOGIC;
                signal internal_out_port_from_the_irq_gen :  STD_LOGIC;
                signal internal_out_port_from_the_portconf_pio :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal internal_out_port_from_the_status_led_pio :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal internal_phasedone_from_the_altpll_0 :  STD_LOGIC;
                signal internal_rTx_Dat_0_from_the_OpenMAC_0 :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal internal_rTx_Dat_1_from_the_OpenMAC_0 :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal internal_rTx_En_0_from_the_OpenMAC_0 :  STD_LOGIC;
                signal internal_rTx_En_1_from_the_OpenMAC_0 :  STD_LOGIC;
                signal internal_sce_from_the_epcs_flash_controller_0 :  STD_LOGIC;
                signal internal_sdo_from_the_epcs_flash_controller_0 :  STD_LOGIC;
                signal internal_select_n_to_the_cfi_flash_0 :  STD_LOGIC;
                signal internal_tri_state_bridge_0_address :  STD_LOGIC_VECTOR (22 DOWNTO 0);
                signal internal_tri_state_bridge_0_readn :  STD_LOGIC;
                signal internal_tri_state_bridge_0_writen :  STD_LOGIC;
                signal internal_zs_addr_from_the_sdram_0 :  STD_LOGIC_VECTOR (11 DOWNTO 0);
                signal internal_zs_ba_from_the_sdram_0 :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal internal_zs_cas_n_from_the_sdram_0 :  STD_LOGIC;
                signal internal_zs_cke_from_the_sdram_0 :  STD_LOGIC;
                signal internal_zs_cs_n_from_the_sdram_0 :  STD_LOGIC;
                signal internal_zs_dqm_from_the_sdram_0 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal internal_zs_ras_n_from_the_sdram_0 :  STD_LOGIC;
                signal internal_zs_we_n_from_the_sdram_0 :  STD_LOGIC;
                signal irq_gen_s1_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal irq_gen_s1_chipselect :  STD_LOGIC;
                signal irq_gen_s1_readdata :  STD_LOGIC;
                signal irq_gen_s1_readdata_from_sa :  STD_LOGIC;
                signal irq_gen_s1_reset_n :  STD_LOGIC;
                signal irq_gen_s1_write_n :  STD_LOGIC;
                signal irq_gen_s1_writedata :  STD_LOGIC;
                signal jtag_uart_0_avalon_jtag_slave_address :  STD_LOGIC;
                signal jtag_uart_0_avalon_jtag_slave_chipselect :  STD_LOGIC;
                signal jtag_uart_0_avalon_jtag_slave_dataavailable :  STD_LOGIC;
                signal jtag_uart_0_avalon_jtag_slave_dataavailable_from_sa :  STD_LOGIC;
                signal jtag_uart_0_avalon_jtag_slave_irq :  STD_LOGIC;
                signal jtag_uart_0_avalon_jtag_slave_irq_from_sa :  STD_LOGIC;
                signal jtag_uart_0_avalon_jtag_slave_read_n :  STD_LOGIC;
                signal jtag_uart_0_avalon_jtag_slave_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal jtag_uart_0_avalon_jtag_slave_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal jtag_uart_0_avalon_jtag_slave_readyfordata :  STD_LOGIC;
                signal jtag_uart_0_avalon_jtag_slave_readyfordata_from_sa :  STD_LOGIC;
                signal jtag_uart_0_avalon_jtag_slave_reset_n :  STD_LOGIC;
                signal jtag_uart_0_avalon_jtag_slave_waitrequest :  STD_LOGIC;
                signal jtag_uart_0_avalon_jtag_slave_waitrequest_from_sa :  STD_LOGIC;
                signal jtag_uart_0_avalon_jtag_slave_write_n :  STD_LOGIC;
                signal jtag_uart_0_avalon_jtag_slave_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal jtag_uart_1_avalon_jtag_slave_address :  STD_LOGIC;
                signal jtag_uart_1_avalon_jtag_slave_chipselect :  STD_LOGIC;
                signal jtag_uart_1_avalon_jtag_slave_dataavailable :  STD_LOGIC;
                signal jtag_uart_1_avalon_jtag_slave_dataavailable_from_sa :  STD_LOGIC;
                signal jtag_uart_1_avalon_jtag_slave_irq :  STD_LOGIC;
                signal jtag_uart_1_avalon_jtag_slave_irq_from_sa :  STD_LOGIC;
                signal jtag_uart_1_avalon_jtag_slave_read_n :  STD_LOGIC;
                signal jtag_uart_1_avalon_jtag_slave_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal jtag_uart_1_avalon_jtag_slave_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal jtag_uart_1_avalon_jtag_slave_readyfordata :  STD_LOGIC;
                signal jtag_uart_1_avalon_jtag_slave_readyfordata_from_sa :  STD_LOGIC;
                signal jtag_uart_1_avalon_jtag_slave_reset_n :  STD_LOGIC;
                signal jtag_uart_1_avalon_jtag_slave_waitrequest :  STD_LOGIC;
                signal jtag_uart_1_avalon_jtag_slave_waitrequest_from_sa :  STD_LOGIC;
                signal jtag_uart_1_avalon_jtag_slave_write_n :  STD_LOGIC;
                signal jtag_uart_1_avalon_jtag_slave_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal module_input12 :  STD_LOGIC;
                signal module_input13 :  STD_LOGIC;
                signal module_input14 :  STD_LOGIC;
                signal module_input15 :  STD_LOGIC;
                signal niosII_openMac_clock_0_in_address :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal niosII_openMac_clock_0_in_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_openMac_clock_0_in_endofpacket :  STD_LOGIC;
                signal niosII_openMac_clock_0_in_endofpacket_from_sa :  STD_LOGIC;
                signal niosII_openMac_clock_0_in_nativeaddress :  STD_LOGIC;
                signal niosII_openMac_clock_0_in_read :  STD_LOGIC;
                signal niosII_openMac_clock_0_in_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal niosII_openMac_clock_0_in_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal niosII_openMac_clock_0_in_reset_n :  STD_LOGIC;
                signal niosII_openMac_clock_0_in_waitrequest :  STD_LOGIC;
                signal niosII_openMac_clock_0_in_waitrequest_from_sa :  STD_LOGIC;
                signal niosII_openMac_clock_0_in_write :  STD_LOGIC;
                signal niosII_openMac_clock_0_in_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal niosII_openMac_clock_0_out_address :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal niosII_openMac_clock_0_out_address_to_slave :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal niosII_openMac_clock_0_out_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_openMac_clock_0_out_endofpacket :  STD_LOGIC;
                signal niosII_openMac_clock_0_out_granted_jtag_uart_0_avalon_jtag_slave :  STD_LOGIC;
                signal niosII_openMac_clock_0_out_nativeaddress :  STD_LOGIC;
                signal niosII_openMac_clock_0_out_qualified_request_jtag_uart_0_avalon_jtag_slave :  STD_LOGIC;
                signal niosII_openMac_clock_0_out_read :  STD_LOGIC;
                signal niosII_openMac_clock_0_out_read_data_valid_jtag_uart_0_avalon_jtag_slave :  STD_LOGIC;
                signal niosII_openMac_clock_0_out_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal niosII_openMac_clock_0_out_requests_jtag_uart_0_avalon_jtag_slave :  STD_LOGIC;
                signal niosII_openMac_clock_0_out_reset_n :  STD_LOGIC;
                signal niosII_openMac_clock_0_out_waitrequest :  STD_LOGIC;
                signal niosII_openMac_clock_0_out_write :  STD_LOGIC;
                signal niosII_openMac_clock_0_out_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal niosII_openMac_clock_1_in_address :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal niosII_openMac_clock_1_in_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_openMac_clock_1_in_endofpacket :  STD_LOGIC;
                signal niosII_openMac_clock_1_in_endofpacket_from_sa :  STD_LOGIC;
                signal niosII_openMac_clock_1_in_nativeaddress :  STD_LOGIC;
                signal niosII_openMac_clock_1_in_read :  STD_LOGIC;
                signal niosII_openMac_clock_1_in_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal niosII_openMac_clock_1_in_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal niosII_openMac_clock_1_in_reset_n :  STD_LOGIC;
                signal niosII_openMac_clock_1_in_waitrequest :  STD_LOGIC;
                signal niosII_openMac_clock_1_in_waitrequest_from_sa :  STD_LOGIC;
                signal niosII_openMac_clock_1_in_write :  STD_LOGIC;
                signal niosII_openMac_clock_1_in_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal niosII_openMac_clock_1_out_address :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal niosII_openMac_clock_1_out_address_to_slave :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal niosII_openMac_clock_1_out_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_openMac_clock_1_out_endofpacket :  STD_LOGIC;
                signal niosII_openMac_clock_1_out_granted_OpenMAC_0_CMP :  STD_LOGIC;
                signal niosII_openMac_clock_1_out_nativeaddress :  STD_LOGIC;
                signal niosII_openMac_clock_1_out_qualified_request_OpenMAC_0_CMP :  STD_LOGIC;
                signal niosII_openMac_clock_1_out_read :  STD_LOGIC;
                signal niosII_openMac_clock_1_out_read_data_valid_OpenMAC_0_CMP :  STD_LOGIC;
                signal niosII_openMac_clock_1_out_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal niosII_openMac_clock_1_out_requests_OpenMAC_0_CMP :  STD_LOGIC;
                signal niosII_openMac_clock_1_out_reset_n :  STD_LOGIC;
                signal niosII_openMac_clock_1_out_waitrequest :  STD_LOGIC;
                signal niosII_openMac_clock_1_out_write :  STD_LOGIC;
                signal niosII_openMac_clock_1_out_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal niosII_openMac_clock_2_in_address :  STD_LOGIC_VECTOR (12 DOWNTO 0);
                signal niosII_openMac_clock_2_in_byteenable :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal niosII_openMac_clock_2_in_endofpacket :  STD_LOGIC;
                signal niosII_openMac_clock_2_in_endofpacket_from_sa :  STD_LOGIC;
                signal niosII_openMac_clock_2_in_nativeaddress :  STD_LOGIC_VECTOR (11 DOWNTO 0);
                signal niosII_openMac_clock_2_in_read :  STD_LOGIC;
                signal niosII_openMac_clock_2_in_readdata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal niosII_openMac_clock_2_in_readdata_from_sa :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal niosII_openMac_clock_2_in_reset_n :  STD_LOGIC;
                signal niosII_openMac_clock_2_in_waitrequest :  STD_LOGIC;
                signal niosII_openMac_clock_2_in_waitrequest_from_sa :  STD_LOGIC;
                signal niosII_openMac_clock_2_in_write :  STD_LOGIC;
                signal niosII_openMac_clock_2_in_writedata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal niosII_openMac_clock_2_out_address :  STD_LOGIC_VECTOR (12 DOWNTO 0);
                signal niosII_openMac_clock_2_out_address_to_slave :  STD_LOGIC_VECTOR (12 DOWNTO 0);
                signal niosII_openMac_clock_2_out_byteenable :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal niosII_openMac_clock_2_out_endofpacket :  STD_LOGIC;
                signal niosII_openMac_clock_2_out_granted_OpenMAC_0_REG :  STD_LOGIC;
                signal niosII_openMac_clock_2_out_nativeaddress :  STD_LOGIC_VECTOR (11 DOWNTO 0);
                signal niosII_openMac_clock_2_out_qualified_request_OpenMAC_0_REG :  STD_LOGIC;
                signal niosII_openMac_clock_2_out_read :  STD_LOGIC;
                signal niosII_openMac_clock_2_out_read_data_valid_OpenMAC_0_REG :  STD_LOGIC;
                signal niosII_openMac_clock_2_out_readdata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal niosII_openMac_clock_2_out_requests_OpenMAC_0_REG :  STD_LOGIC;
                signal niosII_openMac_clock_2_out_reset_n :  STD_LOGIC;
                signal niosII_openMac_clock_2_out_waitrequest :  STD_LOGIC;
                signal niosII_openMac_clock_2_out_write :  STD_LOGIC;
                signal niosII_openMac_clock_2_out_writedata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal niosII_openMac_clock_3_in_address :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_openMac_clock_3_in_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_openMac_clock_3_in_endofpacket :  STD_LOGIC;
                signal niosII_openMac_clock_3_in_endofpacket_from_sa :  STD_LOGIC;
                signal niosII_openMac_clock_3_in_nativeaddress :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal niosII_openMac_clock_3_in_read :  STD_LOGIC;
                signal niosII_openMac_clock_3_in_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal niosII_openMac_clock_3_in_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal niosII_openMac_clock_3_in_reset_n :  STD_LOGIC;
                signal niosII_openMac_clock_3_in_waitrequest :  STD_LOGIC;
                signal niosII_openMac_clock_3_in_waitrequest_from_sa :  STD_LOGIC;
                signal niosII_openMac_clock_3_in_write :  STD_LOGIC;
                signal niosII_openMac_clock_3_in_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal niosII_openMac_clock_3_out_address :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_openMac_clock_3_out_address_to_slave :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_openMac_clock_3_out_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_openMac_clock_3_out_endofpacket :  STD_LOGIC;
                signal niosII_openMac_clock_3_out_granted_altpll_0_pll_slave :  STD_LOGIC;
                signal niosII_openMac_clock_3_out_nativeaddress :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal niosII_openMac_clock_3_out_qualified_request_altpll_0_pll_slave :  STD_LOGIC;
                signal niosII_openMac_clock_3_out_read :  STD_LOGIC;
                signal niosII_openMac_clock_3_out_read_data_valid_altpll_0_pll_slave :  STD_LOGIC;
                signal niosII_openMac_clock_3_out_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal niosII_openMac_clock_3_out_requests_altpll_0_pll_slave :  STD_LOGIC;
                signal niosII_openMac_clock_3_out_reset_n :  STD_LOGIC;
                signal niosII_openMac_clock_3_out_waitrequest :  STD_LOGIC;
                signal niosII_openMac_clock_3_out_write :  STD_LOGIC;
                signal niosII_openMac_clock_3_out_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal niosII_openMac_clock_4_in_address :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal niosII_openMac_clock_4_in_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_openMac_clock_4_in_endofpacket :  STD_LOGIC;
                signal niosII_openMac_clock_4_in_endofpacket_from_sa :  STD_LOGIC;
                signal niosII_openMac_clock_4_in_nativeaddress :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal niosII_openMac_clock_4_in_read :  STD_LOGIC;
                signal niosII_openMac_clock_4_in_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal niosII_openMac_clock_4_in_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal niosII_openMac_clock_4_in_reset_n :  STD_LOGIC;
                signal niosII_openMac_clock_4_in_waitrequest :  STD_LOGIC;
                signal niosII_openMac_clock_4_in_waitrequest_from_sa :  STD_LOGIC;
                signal niosII_openMac_clock_4_in_write :  STD_LOGIC;
                signal niosII_openMac_clock_4_in_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal niosII_openMac_clock_4_out_address :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal niosII_openMac_clock_4_out_address_to_slave :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal niosII_openMac_clock_4_out_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal niosII_openMac_clock_4_out_endofpacket :  STD_LOGIC;
                signal niosII_openMac_clock_4_out_granted_remote_update_cycloneiii_0_s1 :  STD_LOGIC;
                signal niosII_openMac_clock_4_out_nativeaddress :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal niosII_openMac_clock_4_out_qualified_request_remote_update_cycloneiii_0_s1 :  STD_LOGIC;
                signal niosII_openMac_clock_4_out_read :  STD_LOGIC;
                signal niosII_openMac_clock_4_out_read_data_valid_remote_update_cycloneiii_0_s1 :  STD_LOGIC;
                signal niosII_openMac_clock_4_out_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal niosII_openMac_clock_4_out_requests_remote_update_cycloneiii_0_s1 :  STD_LOGIC;
                signal niosII_openMac_clock_4_out_reset_n :  STD_LOGIC;
                signal niosII_openMac_clock_4_out_waitrequest :  STD_LOGIC;
                signal niosII_openMac_clock_4_out_write :  STD_LOGIC;
                signal niosII_openMac_clock_4_out_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal node_switch_pio_s1_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal node_switch_pio_s1_readdata :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal node_switch_pio_s1_readdata_from_sa :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal node_switch_pio_s1_reset_n :  STD_LOGIC;
                signal onchip_memory_0_s1_address :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal onchip_memory_0_s1_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal onchip_memory_0_s1_chipselect :  STD_LOGIC;
                signal onchip_memory_0_s1_clken :  STD_LOGIC;
                signal onchip_memory_0_s1_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal onchip_memory_0_s1_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal onchip_memory_0_s1_write :  STD_LOGIC;
                signal onchip_memory_0_s1_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal out_clk_altpll_0_c0 :  STD_LOGIC;
                signal out_clk_altpll_0_c1 :  STD_LOGIC;
                signal out_clk_altpll_0_c2 :  STD_LOGIC;
                signal out_clk_altpll_0_c3 :  STD_LOGIC;
                signal out_clk_altpll_0_c4 :  STD_LOGIC;
                signal pcp_cpu_data_master_address :  STD_LOGIC_VECTOR (25 DOWNTO 0);
                signal pcp_cpu_data_master_address_to_slave :  STD_LOGIC_VECTOR (25 DOWNTO 0);
                signal pcp_cpu_data_master_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal pcp_cpu_data_master_byteenable_DBC3C40_SRAM_0_avalon_tristate_slave :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal pcp_cpu_data_master_byteenable_cfi_flash_0_s1 :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal pcp_cpu_data_master_byteenable_niosII_openMac_clock_2_in :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal pcp_cpu_data_master_dbs_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal pcp_cpu_data_master_dbs_write_16 :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal pcp_cpu_data_master_debugaccess :  STD_LOGIC;
                signal pcp_cpu_data_master_granted_DBC3C40_SRAM_0_avalon_tristate_slave :  STD_LOGIC;
                signal pcp_cpu_data_master_granted_OpenMAC_0_iBuf :  STD_LOGIC;
                signal pcp_cpu_data_master_granted_cfi_flash_0_s1 :  STD_LOGIC;
                signal pcp_cpu_data_master_granted_clock_crossing_0_s1 :  STD_LOGIC;
                signal pcp_cpu_data_master_granted_cnApi_Av2Av_0_pcp :  STD_LOGIC;
                signal pcp_cpu_data_master_granted_epcs_flash_controller_0_epcs_control_port :  STD_LOGIC;
                signal pcp_cpu_data_master_granted_niosII_openMac_clock_0_in :  STD_LOGIC;
                signal pcp_cpu_data_master_granted_niosII_openMac_clock_1_in :  STD_LOGIC;
                signal pcp_cpu_data_master_granted_niosII_openMac_clock_2_in :  STD_LOGIC;
                signal pcp_cpu_data_master_granted_niosII_openMac_clock_3_in :  STD_LOGIC;
                signal pcp_cpu_data_master_granted_niosII_openMac_clock_4_in :  STD_LOGIC;
                signal pcp_cpu_data_master_granted_onchip_memory_0_s1 :  STD_LOGIC;
                signal pcp_cpu_data_master_granted_pcp_cpu_jtag_debug_module :  STD_LOGIC;
                signal pcp_cpu_data_master_irq :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal pcp_cpu_data_master_no_byte_enables_and_last_term :  STD_LOGIC;
                signal pcp_cpu_data_master_qualified_request_DBC3C40_SRAM_0_avalon_tristate_slave :  STD_LOGIC;
                signal pcp_cpu_data_master_qualified_request_OpenMAC_0_iBuf :  STD_LOGIC;
                signal pcp_cpu_data_master_qualified_request_cfi_flash_0_s1 :  STD_LOGIC;
                signal pcp_cpu_data_master_qualified_request_clock_crossing_0_s1 :  STD_LOGIC;
                signal pcp_cpu_data_master_qualified_request_cnApi_Av2Av_0_pcp :  STD_LOGIC;
                signal pcp_cpu_data_master_qualified_request_epcs_flash_controller_0_epcs_control_port :  STD_LOGIC;
                signal pcp_cpu_data_master_qualified_request_niosII_openMac_clock_0_in :  STD_LOGIC;
                signal pcp_cpu_data_master_qualified_request_niosII_openMac_clock_1_in :  STD_LOGIC;
                signal pcp_cpu_data_master_qualified_request_niosII_openMac_clock_2_in :  STD_LOGIC;
                signal pcp_cpu_data_master_qualified_request_niosII_openMac_clock_3_in :  STD_LOGIC;
                signal pcp_cpu_data_master_qualified_request_niosII_openMac_clock_4_in :  STD_LOGIC;
                signal pcp_cpu_data_master_qualified_request_onchip_memory_0_s1 :  STD_LOGIC;
                signal pcp_cpu_data_master_qualified_request_pcp_cpu_jtag_debug_module :  STD_LOGIC;
                signal pcp_cpu_data_master_read :  STD_LOGIC;
                signal pcp_cpu_data_master_read_data_valid_DBC3C40_SRAM_0_avalon_tristate_slave :  STD_LOGIC;
                signal pcp_cpu_data_master_read_data_valid_OpenMAC_0_iBuf :  STD_LOGIC;
                signal pcp_cpu_data_master_read_data_valid_cfi_flash_0_s1 :  STD_LOGIC;
                signal pcp_cpu_data_master_read_data_valid_clock_crossing_0_s1 :  STD_LOGIC;
                signal pcp_cpu_data_master_read_data_valid_clock_crossing_0_s1_shift_register :  STD_LOGIC;
                signal pcp_cpu_data_master_read_data_valid_cnApi_Av2Av_0_pcp :  STD_LOGIC;
                signal pcp_cpu_data_master_read_data_valid_epcs_flash_controller_0_epcs_control_port :  STD_LOGIC;
                signal pcp_cpu_data_master_read_data_valid_niosII_openMac_clock_0_in :  STD_LOGIC;
                signal pcp_cpu_data_master_read_data_valid_niosII_openMac_clock_1_in :  STD_LOGIC;
                signal pcp_cpu_data_master_read_data_valid_niosII_openMac_clock_2_in :  STD_LOGIC;
                signal pcp_cpu_data_master_read_data_valid_niosII_openMac_clock_3_in :  STD_LOGIC;
                signal pcp_cpu_data_master_read_data_valid_niosII_openMac_clock_4_in :  STD_LOGIC;
                signal pcp_cpu_data_master_read_data_valid_onchip_memory_0_s1 :  STD_LOGIC;
                signal pcp_cpu_data_master_read_data_valid_pcp_cpu_jtag_debug_module :  STD_LOGIC;
                signal pcp_cpu_data_master_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal pcp_cpu_data_master_requests_DBC3C40_SRAM_0_avalon_tristate_slave :  STD_LOGIC;
                signal pcp_cpu_data_master_requests_OpenMAC_0_iBuf :  STD_LOGIC;
                signal pcp_cpu_data_master_requests_cfi_flash_0_s1 :  STD_LOGIC;
                signal pcp_cpu_data_master_requests_clock_crossing_0_s1 :  STD_LOGIC;
                signal pcp_cpu_data_master_requests_cnApi_Av2Av_0_pcp :  STD_LOGIC;
                signal pcp_cpu_data_master_requests_epcs_flash_controller_0_epcs_control_port :  STD_LOGIC;
                signal pcp_cpu_data_master_requests_niosII_openMac_clock_0_in :  STD_LOGIC;
                signal pcp_cpu_data_master_requests_niosII_openMac_clock_1_in :  STD_LOGIC;
                signal pcp_cpu_data_master_requests_niosII_openMac_clock_2_in :  STD_LOGIC;
                signal pcp_cpu_data_master_requests_niosII_openMac_clock_3_in :  STD_LOGIC;
                signal pcp_cpu_data_master_requests_niosII_openMac_clock_4_in :  STD_LOGIC;
                signal pcp_cpu_data_master_requests_onchip_memory_0_s1 :  STD_LOGIC;
                signal pcp_cpu_data_master_requests_pcp_cpu_jtag_debug_module :  STD_LOGIC;
                signal pcp_cpu_data_master_waitrequest :  STD_LOGIC;
                signal pcp_cpu_data_master_write :  STD_LOGIC;
                signal pcp_cpu_data_master_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal pcp_cpu_instruction_master_address :  STD_LOGIC_VECTOR (25 DOWNTO 0);
                signal pcp_cpu_instruction_master_address_to_slave :  STD_LOGIC_VECTOR (25 DOWNTO 0);
                signal pcp_cpu_instruction_master_dbs_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal pcp_cpu_instruction_master_granted_DBC3C40_SRAM_0_avalon_tristate_slave :  STD_LOGIC;
                signal pcp_cpu_instruction_master_granted_cfi_flash_0_s1 :  STD_LOGIC;
                signal pcp_cpu_instruction_master_granted_epcs_flash_controller_0_epcs_control_port :  STD_LOGIC;
                signal pcp_cpu_instruction_master_granted_onchip_memory_0_s1 :  STD_LOGIC;
                signal pcp_cpu_instruction_master_granted_pcp_cpu_jtag_debug_module :  STD_LOGIC;
                signal pcp_cpu_instruction_master_latency_counter :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal pcp_cpu_instruction_master_qualified_request_DBC3C40_SRAM_0_avalon_tristate_slave :  STD_LOGIC;
                signal pcp_cpu_instruction_master_qualified_request_cfi_flash_0_s1 :  STD_LOGIC;
                signal pcp_cpu_instruction_master_qualified_request_epcs_flash_controller_0_epcs_control_port :  STD_LOGIC;
                signal pcp_cpu_instruction_master_qualified_request_onchip_memory_0_s1 :  STD_LOGIC;
                signal pcp_cpu_instruction_master_qualified_request_pcp_cpu_jtag_debug_module :  STD_LOGIC;
                signal pcp_cpu_instruction_master_read :  STD_LOGIC;
                signal pcp_cpu_instruction_master_read_data_valid_DBC3C40_SRAM_0_avalon_tristate_slave :  STD_LOGIC;
                signal pcp_cpu_instruction_master_read_data_valid_cfi_flash_0_s1 :  STD_LOGIC;
                signal pcp_cpu_instruction_master_read_data_valid_epcs_flash_controller_0_epcs_control_port :  STD_LOGIC;
                signal pcp_cpu_instruction_master_read_data_valid_onchip_memory_0_s1 :  STD_LOGIC;
                signal pcp_cpu_instruction_master_read_data_valid_pcp_cpu_jtag_debug_module :  STD_LOGIC;
                signal pcp_cpu_instruction_master_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal pcp_cpu_instruction_master_readdatavalid :  STD_LOGIC;
                signal pcp_cpu_instruction_master_requests_DBC3C40_SRAM_0_avalon_tristate_slave :  STD_LOGIC;
                signal pcp_cpu_instruction_master_requests_cfi_flash_0_s1 :  STD_LOGIC;
                signal pcp_cpu_instruction_master_requests_epcs_flash_controller_0_epcs_control_port :  STD_LOGIC;
                signal pcp_cpu_instruction_master_requests_onchip_memory_0_s1 :  STD_LOGIC;
                signal pcp_cpu_instruction_master_requests_pcp_cpu_jtag_debug_module :  STD_LOGIC;
                signal pcp_cpu_instruction_master_waitrequest :  STD_LOGIC;
                signal pcp_cpu_jtag_debug_module_address :  STD_LOGIC_VECTOR (8 DOWNTO 0);
                signal pcp_cpu_jtag_debug_module_begintransfer :  STD_LOGIC;
                signal pcp_cpu_jtag_debug_module_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal pcp_cpu_jtag_debug_module_chipselect :  STD_LOGIC;
                signal pcp_cpu_jtag_debug_module_debugaccess :  STD_LOGIC;
                signal pcp_cpu_jtag_debug_module_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal pcp_cpu_jtag_debug_module_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal pcp_cpu_jtag_debug_module_reset_n :  STD_LOGIC;
                signal pcp_cpu_jtag_debug_module_resetrequest :  STD_LOGIC;
                signal pcp_cpu_jtag_debug_module_resetrequest_from_sa :  STD_LOGIC;
                signal pcp_cpu_jtag_debug_module_write :  STD_LOGIC;
                signal pcp_cpu_jtag_debug_module_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal portconf_pio_s1_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal portconf_pio_s1_chipselect :  STD_LOGIC;
                signal portconf_pio_s1_readdata :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal portconf_pio_s1_readdata_from_sa :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal portconf_pio_s1_reset_n :  STD_LOGIC;
                signal portconf_pio_s1_write_n :  STD_LOGIC;
                signal portconf_pio_s1_writedata :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal registered_pcp_cpu_data_master_read_data_valid_DBC3C40_SRAM_0_avalon_tristate_slave :  STD_LOGIC;
                signal registered_pcp_cpu_data_master_read_data_valid_cfi_flash_0_s1 :  STD_LOGIC;
                signal registered_pcp_cpu_data_master_read_data_valid_onchip_memory_0_s1 :  STD_LOGIC;
                signal remote_update_cycloneiii_0_s1_address :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal remote_update_cycloneiii_0_s1_chipselect :  STD_LOGIC;
                signal remote_update_cycloneiii_0_s1_read :  STD_LOGIC;
                signal remote_update_cycloneiii_0_s1_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal remote_update_cycloneiii_0_s1_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal remote_update_cycloneiii_0_s1_reset :  STD_LOGIC;
                signal remote_update_cycloneiii_0_s1_waitrequest :  STD_LOGIC;
                signal remote_update_cycloneiii_0_s1_waitrequest_from_sa :  STD_LOGIC;
                signal remote_update_cycloneiii_0_s1_write :  STD_LOGIC;
                signal remote_update_cycloneiii_0_s1_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal reset_n_sources :  STD_LOGIC;
                signal sdram_0_s1_address :  STD_LOGIC_VECTOR (21 DOWNTO 0);
                signal sdram_0_s1_byteenable_n :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal sdram_0_s1_chipselect :  STD_LOGIC;
                signal sdram_0_s1_read_n :  STD_LOGIC;
                signal sdram_0_s1_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal sdram_0_s1_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal sdram_0_s1_readdatavalid :  STD_LOGIC;
                signal sdram_0_s1_reset_n :  STD_LOGIC;
                signal sdram_0_s1_waitrequest :  STD_LOGIC;
                signal sdram_0_s1_waitrequest_from_sa :  STD_LOGIC;
                signal sdram_0_s1_write_n :  STD_LOGIC;
                signal sdram_0_s1_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal status_led_pio_s1_address :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal status_led_pio_s1_chipselect :  STD_LOGIC;
                signal status_led_pio_s1_readdata :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal status_led_pio_s1_readdata_from_sa :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal status_led_pio_s1_reset_n :  STD_LOGIC;
                signal status_led_pio_s1_write_n :  STD_LOGIC;
                signal status_led_pio_s1_writedata :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal sync_irq_s1_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal sync_irq_s1_chipselect :  STD_LOGIC;
                signal sync_irq_s1_irq :  STD_LOGIC;
                signal sync_irq_s1_irq_from_sa :  STD_LOGIC;
                signal sync_irq_s1_readdata :  STD_LOGIC;
                signal sync_irq_s1_readdata_from_sa :  STD_LOGIC;
                signal sync_irq_s1_reset_n :  STD_LOGIC;
                signal sync_irq_s1_write_n :  STD_LOGIC;
                signal sync_irq_s1_writedata :  STD_LOGIC;
                signal sysid_control_slave_address :  STD_LOGIC;
                signal sysid_control_slave_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal sysid_control_slave_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal system_timer_ap_s1_address :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal system_timer_ap_s1_chipselect :  STD_LOGIC;
                signal system_timer_ap_s1_irq :  STD_LOGIC;
                signal system_timer_ap_s1_irq_from_sa :  STD_LOGIC;
                signal system_timer_ap_s1_readdata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal system_timer_ap_s1_readdata_from_sa :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal system_timer_ap_s1_reset_n :  STD_LOGIC;
                signal system_timer_ap_s1_write_n :  STD_LOGIC;
                signal system_timer_ap_s1_writedata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal system_timer_s1_address :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal system_timer_s1_chipselect :  STD_LOGIC;
                signal system_timer_s1_irq :  STD_LOGIC;
                signal system_timer_s1_irq_from_sa :  STD_LOGIC;
                signal system_timer_s1_readdata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal system_timer_s1_readdata_from_sa :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal system_timer_s1_reset_n :  STD_LOGIC;
                signal system_timer_s1_write_n :  STD_LOGIC;
                signal system_timer_s1_writedata :  STD_LOGIC_VECTOR (15 DOWNTO 0);

begin

  --the_OpenMAC_0_CMP, which is an e_instance
  the_OpenMAC_0_CMP : OpenMAC_0_CMP_arbitrator
    port map(
      OpenMAC_0_CMP_address => OpenMAC_0_CMP_address,
      OpenMAC_0_CMP_byteenable_n => OpenMAC_0_CMP_byteenable_n,
      OpenMAC_0_CMP_chipselect => OpenMAC_0_CMP_chipselect,
      OpenMAC_0_CMP_irq_from_sa => OpenMAC_0_CMP_irq_from_sa,
      OpenMAC_0_CMP_read_n => OpenMAC_0_CMP_read_n,
      OpenMAC_0_CMP_readdata_from_sa => OpenMAC_0_CMP_readdata_from_sa,
      OpenMAC_0_CMP_reset_n => OpenMAC_0_CMP_reset_n,
      OpenMAC_0_CMP_write_n => OpenMAC_0_CMP_write_n,
      OpenMAC_0_CMP_writedata => OpenMAC_0_CMP_writedata,
      d1_OpenMAC_0_CMP_end_xfer => d1_OpenMAC_0_CMP_end_xfer,
      niosII_openMac_clock_1_out_granted_OpenMAC_0_CMP => niosII_openMac_clock_1_out_granted_OpenMAC_0_CMP,
      niosII_openMac_clock_1_out_qualified_request_OpenMAC_0_CMP => niosII_openMac_clock_1_out_qualified_request_OpenMAC_0_CMP,
      niosII_openMac_clock_1_out_read_data_valid_OpenMAC_0_CMP => niosII_openMac_clock_1_out_read_data_valid_OpenMAC_0_CMP,
      niosII_openMac_clock_1_out_requests_OpenMAC_0_CMP => niosII_openMac_clock_1_out_requests_OpenMAC_0_CMP,
      OpenMAC_0_CMP_irq => OpenMAC_0_CMP_irq,
      OpenMAC_0_CMP_readdata => OpenMAC_0_CMP_readdata,
      clk => internal_clk50Meg,
      niosII_openMac_clock_1_out_address_to_slave => niosII_openMac_clock_1_out_address_to_slave,
      niosII_openMac_clock_1_out_byteenable => niosII_openMac_clock_1_out_byteenable,
      niosII_openMac_clock_1_out_read => niosII_openMac_clock_1_out_read,
      niosII_openMac_clock_1_out_write => niosII_openMac_clock_1_out_write,
      niosII_openMac_clock_1_out_writedata => niosII_openMac_clock_1_out_writedata,
      reset_n => clk50Meg_reset_n
    );


  --the_OpenMAC_0_REG, which is an e_instance
  the_OpenMAC_0_REG : OpenMAC_0_REG_arbitrator
    port map(
      OpenMAC_0_REG_address => OpenMAC_0_REG_address,
      OpenMAC_0_REG_byteenable_n => OpenMAC_0_REG_byteenable_n,
      OpenMAC_0_REG_chipselect => OpenMAC_0_REG_chipselect,
      OpenMAC_0_REG_irq_from_sa => OpenMAC_0_REG_irq_from_sa,
      OpenMAC_0_REG_read_n => OpenMAC_0_REG_read_n,
      OpenMAC_0_REG_readdata_from_sa => OpenMAC_0_REG_readdata_from_sa,
      OpenMAC_0_REG_write_n => OpenMAC_0_REG_write_n,
      OpenMAC_0_REG_writedata => OpenMAC_0_REG_writedata,
      d1_OpenMAC_0_REG_end_xfer => d1_OpenMAC_0_REG_end_xfer,
      niosII_openMac_clock_2_out_granted_OpenMAC_0_REG => niosII_openMac_clock_2_out_granted_OpenMAC_0_REG,
      niosII_openMac_clock_2_out_qualified_request_OpenMAC_0_REG => niosII_openMac_clock_2_out_qualified_request_OpenMAC_0_REG,
      niosII_openMac_clock_2_out_read_data_valid_OpenMAC_0_REG => niosII_openMac_clock_2_out_read_data_valid_OpenMAC_0_REG,
      niosII_openMac_clock_2_out_requests_OpenMAC_0_REG => niosII_openMac_clock_2_out_requests_OpenMAC_0_REG,
      OpenMAC_0_REG_irq => OpenMAC_0_REG_irq,
      OpenMAC_0_REG_readdata => OpenMAC_0_REG_readdata,
      clk => internal_clk50Meg,
      niosII_openMac_clock_2_out_address_to_slave => niosII_openMac_clock_2_out_address_to_slave,
      niosII_openMac_clock_2_out_byteenable => niosII_openMac_clock_2_out_byteenable,
      niosII_openMac_clock_2_out_read => niosII_openMac_clock_2_out_read,
      niosII_openMac_clock_2_out_write => niosII_openMac_clock_2_out_write,
      niosII_openMac_clock_2_out_writedata => niosII_openMac_clock_2_out_writedata,
      reset_n => clk50Meg_reset_n
    );


  --the_OpenMAC_0_iBuf, which is an e_instance
  the_OpenMAC_0_iBuf : OpenMAC_0_iBuf_arbitrator
    port map(
      OpenMAC_0_iBuf_address => OpenMAC_0_iBuf_address,
      OpenMAC_0_iBuf_byteenable => OpenMAC_0_iBuf_byteenable,
      OpenMAC_0_iBuf_chipselect => OpenMAC_0_iBuf_chipselect,
      OpenMAC_0_iBuf_read_n => OpenMAC_0_iBuf_read_n,
      OpenMAC_0_iBuf_readdata_from_sa => OpenMAC_0_iBuf_readdata_from_sa,
      OpenMAC_0_iBuf_wait_counter_eq_0 => OpenMAC_0_iBuf_wait_counter_eq_0,
      OpenMAC_0_iBuf_write_n => OpenMAC_0_iBuf_write_n,
      OpenMAC_0_iBuf_writedata => OpenMAC_0_iBuf_writedata,
      d1_OpenMAC_0_iBuf_end_xfer => d1_OpenMAC_0_iBuf_end_xfer,
      pcp_cpu_data_master_granted_OpenMAC_0_iBuf => pcp_cpu_data_master_granted_OpenMAC_0_iBuf,
      pcp_cpu_data_master_qualified_request_OpenMAC_0_iBuf => pcp_cpu_data_master_qualified_request_OpenMAC_0_iBuf,
      pcp_cpu_data_master_read_data_valid_OpenMAC_0_iBuf => pcp_cpu_data_master_read_data_valid_OpenMAC_0_iBuf,
      pcp_cpu_data_master_requests_OpenMAC_0_iBuf => pcp_cpu_data_master_requests_OpenMAC_0_iBuf,
      OpenMAC_0_iBuf_readdata => OpenMAC_0_iBuf_readdata,
      clk => internal_clk90Meg,
      pcp_cpu_data_master_address_to_slave => pcp_cpu_data_master_address_to_slave,
      pcp_cpu_data_master_byteenable => pcp_cpu_data_master_byteenable,
      pcp_cpu_data_master_read => pcp_cpu_data_master_read,
      pcp_cpu_data_master_waitrequest => pcp_cpu_data_master_waitrequest,
      pcp_cpu_data_master_write => pcp_cpu_data_master_write,
      pcp_cpu_data_master_writedata => pcp_cpu_data_master_writedata,
      reset_n => clk90Meg_reset_n
    );


  --the_OpenMAC_0, which is an e_ptf_instance
  the_OpenMAC_0 : OpenMAC_0
    port map(
      iBuf_readdata => OpenMAC_0_iBuf_readdata,
      mii_Clk => internal_mii_Clk_from_the_OpenMAC_0,
      mii_Do => internal_mii_Do_from_the_OpenMAC_0,
      mii_Doe => internal_mii_Doe_from_the_OpenMAC_0,
      mii_nResetOut => internal_mii_nResetOut_from_the_OpenMAC_0,
      rTx_Dat_0 => internal_rTx_Dat_0_from_the_OpenMAC_0,
      rTx_Dat_1 => internal_rTx_Dat_1_from_the_OpenMAC_0,
      rTx_En_0 => internal_rTx_En_0_from_the_OpenMAC_0,
      rTx_En_1 => internal_rTx_En_1_from_the_OpenMAC_0,
      s_IRQ => OpenMAC_0_REG_irq,
      s_readdata => OpenMAC_0_REG_readdata,
      t_IRQ => OpenMAC_0_CMP_irq,
      t_readdata => OpenMAC_0_CMP_readdata,
      Clk50 => internal_clk50Meg,
      ClkFaster => internal_clk90Meg,
      Reset_n => OpenMAC_0_CMP_reset_n,
      iBuf_address => OpenMAC_0_iBuf_address,
      iBuf_byteenable => OpenMAC_0_iBuf_byteenable,
      iBuf_chipselect => OpenMAC_0_iBuf_chipselect,
      iBuf_read_n => OpenMAC_0_iBuf_read_n,
      iBuf_write_n => OpenMAC_0_iBuf_write_n,
      iBuf_writedata => OpenMAC_0_iBuf_writedata,
      mii_Di => mii_Di_to_the_OpenMAC_0,
      rCrs_Dv_0 => rCrs_Dv_0_to_the_OpenMAC_0,
      rCrs_Dv_1 => rCrs_Dv_1_to_the_OpenMAC_0,
      rRx_Dat_0 => rRx_Dat_0_to_the_OpenMAC_0,
      rRx_Dat_1 => rRx_Dat_1_to_the_OpenMAC_0,
      s_address => OpenMAC_0_REG_address,
      s_byteenable_n => OpenMAC_0_REG_byteenable_n,
      s_chipselect => OpenMAC_0_REG_chipselect,
      s_read_n => OpenMAC_0_REG_read_n,
      s_write_n => OpenMAC_0_REG_write_n,
      s_writedata => OpenMAC_0_REG_writedata,
      t_address(0) => OpenMAC_0_CMP_address,
      t_byteenable_n => OpenMAC_0_CMP_byteenable_n,
      t_chipselect => OpenMAC_0_CMP_chipselect,
      t_read_n => OpenMAC_0_CMP_read_n,
      t_write_n => OpenMAC_0_CMP_write_n,
      t_writedata => OpenMAC_0_CMP_writedata
    );


  --the_altpll_0_pll_slave, which is an e_instance
  the_altpll_0_pll_slave : altpll_0_pll_slave_arbitrator
    port map(
      altpll_0_pll_slave_address => altpll_0_pll_slave_address,
      altpll_0_pll_slave_read => altpll_0_pll_slave_read,
      altpll_0_pll_slave_readdata_from_sa => altpll_0_pll_slave_readdata_from_sa,
      altpll_0_pll_slave_reset => altpll_0_pll_slave_reset,
      altpll_0_pll_slave_write => altpll_0_pll_slave_write,
      altpll_0_pll_slave_writedata => altpll_0_pll_slave_writedata,
      d1_altpll_0_pll_slave_end_xfer => d1_altpll_0_pll_slave_end_xfer,
      niosII_openMac_clock_3_out_granted_altpll_0_pll_slave => niosII_openMac_clock_3_out_granted_altpll_0_pll_slave,
      niosII_openMac_clock_3_out_qualified_request_altpll_0_pll_slave => niosII_openMac_clock_3_out_qualified_request_altpll_0_pll_slave,
      niosII_openMac_clock_3_out_read_data_valid_altpll_0_pll_slave => niosII_openMac_clock_3_out_read_data_valid_altpll_0_pll_slave,
      niosII_openMac_clock_3_out_requests_altpll_0_pll_slave => niosII_openMac_clock_3_out_requests_altpll_0_pll_slave,
      altpll_0_pll_slave_readdata => altpll_0_pll_slave_readdata,
      clk => clk_0,
      niosII_openMac_clock_3_out_address_to_slave => niosII_openMac_clock_3_out_address_to_slave,
      niosII_openMac_clock_3_out_read => niosII_openMac_clock_3_out_read,
      niosII_openMac_clock_3_out_write => niosII_openMac_clock_3_out_write,
      niosII_openMac_clock_3_out_writedata => niosII_openMac_clock_3_out_writedata,
      reset_n => clk_0_reset_n
    );


  --clk50Meg out_clk assignment, which is an e_assign
  internal_clk50Meg <= out_clk_altpll_0_c0;
  --clk90Meg out_clk assignment, which is an e_assign
  internal_clk90Meg <= out_clk_altpll_0_c1;
  --clk100Meg180 out_clk assignment, which is an e_assign
  clk100Meg180 <= out_clk_altpll_0_c2;
  --clk90MegSDRAM out_clk assignment, which is an e_assign
  clk90MegSDRAM <= out_clk_altpll_0_c3;
  --clk25Meg out_clk assignment, which is an e_assign
  internal_clk25Meg <= out_clk_altpll_0_c4;
  --the_altpll_0, which is an e_ptf_instance
  the_altpll_0 : altpll_0
    port map(
      c0 => out_clk_altpll_0_c0,
      c1 => out_clk_altpll_0_c1,
      c2 => out_clk_altpll_0_c2,
      c3 => out_clk_altpll_0_c3,
      c4 => out_clk_altpll_0_c4,
      locked => internal_locked_from_the_altpll_0,
      phasedone => internal_phasedone_from_the_altpll_0,
      readdata => altpll_0_pll_slave_readdata,
      address => altpll_0_pll_slave_address,
      clk => clk_0,
      read => altpll_0_pll_slave_read,
      reset => altpll_0_pll_slave_reset,
      write => altpll_0_pll_slave_write,
      writedata => altpll_0_pll_slave_writedata
    );


  --the_ap_cpu_jtag_debug_module, which is an e_instance
  the_ap_cpu_jtag_debug_module : ap_cpu_jtag_debug_module_arbitrator
    port map(
      ap_cpu_data_master_granted_ap_cpu_jtag_debug_module => ap_cpu_data_master_granted_ap_cpu_jtag_debug_module,
      ap_cpu_data_master_qualified_request_ap_cpu_jtag_debug_module => ap_cpu_data_master_qualified_request_ap_cpu_jtag_debug_module,
      ap_cpu_data_master_read_data_valid_ap_cpu_jtag_debug_module => ap_cpu_data_master_read_data_valid_ap_cpu_jtag_debug_module,
      ap_cpu_data_master_requests_ap_cpu_jtag_debug_module => ap_cpu_data_master_requests_ap_cpu_jtag_debug_module,
      ap_cpu_instruction_master_granted_ap_cpu_jtag_debug_module => ap_cpu_instruction_master_granted_ap_cpu_jtag_debug_module,
      ap_cpu_instruction_master_qualified_request_ap_cpu_jtag_debug_module => ap_cpu_instruction_master_qualified_request_ap_cpu_jtag_debug_module,
      ap_cpu_instruction_master_read_data_valid_ap_cpu_jtag_debug_module => ap_cpu_instruction_master_read_data_valid_ap_cpu_jtag_debug_module,
      ap_cpu_instruction_master_requests_ap_cpu_jtag_debug_module => ap_cpu_instruction_master_requests_ap_cpu_jtag_debug_module,
      ap_cpu_jtag_debug_module_address => ap_cpu_jtag_debug_module_address,
      ap_cpu_jtag_debug_module_begintransfer => ap_cpu_jtag_debug_module_begintransfer,
      ap_cpu_jtag_debug_module_byteenable => ap_cpu_jtag_debug_module_byteenable,
      ap_cpu_jtag_debug_module_chipselect => ap_cpu_jtag_debug_module_chipselect,
      ap_cpu_jtag_debug_module_debugaccess => ap_cpu_jtag_debug_module_debugaccess,
      ap_cpu_jtag_debug_module_readdata_from_sa => ap_cpu_jtag_debug_module_readdata_from_sa,
      ap_cpu_jtag_debug_module_reset_n => ap_cpu_jtag_debug_module_reset_n,
      ap_cpu_jtag_debug_module_resetrequest_from_sa => ap_cpu_jtag_debug_module_resetrequest_from_sa,
      ap_cpu_jtag_debug_module_write => ap_cpu_jtag_debug_module_write,
      ap_cpu_jtag_debug_module_writedata => ap_cpu_jtag_debug_module_writedata,
      d1_ap_cpu_jtag_debug_module_end_xfer => d1_ap_cpu_jtag_debug_module_end_xfer,
      ap_cpu_data_master_address_to_slave => ap_cpu_data_master_address_to_slave,
      ap_cpu_data_master_byteenable => ap_cpu_data_master_byteenable,
      ap_cpu_data_master_debugaccess => ap_cpu_data_master_debugaccess,
      ap_cpu_data_master_read => ap_cpu_data_master_read,
      ap_cpu_data_master_waitrequest => ap_cpu_data_master_waitrequest,
      ap_cpu_data_master_write => ap_cpu_data_master_write,
      ap_cpu_data_master_writedata => ap_cpu_data_master_writedata,
      ap_cpu_instruction_master_address_to_slave => ap_cpu_instruction_master_address_to_slave,
      ap_cpu_instruction_master_latency_counter => ap_cpu_instruction_master_latency_counter,
      ap_cpu_instruction_master_read => ap_cpu_instruction_master_read,
      ap_cpu_instruction_master_read_data_valid_sdram_0_s1_shift_register => ap_cpu_instruction_master_read_data_valid_sdram_0_s1_shift_register,
      ap_cpu_jtag_debug_module_readdata => ap_cpu_jtag_debug_module_readdata,
      ap_cpu_jtag_debug_module_resetrequest => ap_cpu_jtag_debug_module_resetrequest,
      clk => internal_clk90Meg,
      reset_n => clk90Meg_reset_n
    );


  --the_ap_cpu_data_master, which is an e_instance
  the_ap_cpu_data_master : ap_cpu_data_master_arbitrator
    port map(
      ap_cpu_data_master_address_to_slave => ap_cpu_data_master_address_to_slave,
      ap_cpu_data_master_irq => ap_cpu_data_master_irq,
      ap_cpu_data_master_readdata => ap_cpu_data_master_readdata,
      ap_cpu_data_master_waitrequest => ap_cpu_data_master_waitrequest,
      ap_cpu_data_master_address => ap_cpu_data_master_address,
      ap_cpu_data_master_granted_ap_cpu_jtag_debug_module => ap_cpu_data_master_granted_ap_cpu_jtag_debug_module,
      ap_cpu_data_master_granted_clock_crossing_1_s1 => ap_cpu_data_master_granted_clock_crossing_1_s1,
      ap_cpu_data_master_granted_cnApi_Av2Av_0_ap => ap_cpu_data_master_granted_cnApi_Av2Av_0_ap,
      ap_cpu_data_master_granted_jtag_uart_1_avalon_jtag_slave => ap_cpu_data_master_granted_jtag_uart_1_avalon_jtag_slave,
      ap_cpu_data_master_granted_sdram_0_s1 => ap_cpu_data_master_granted_sdram_0_s1,
      ap_cpu_data_master_qualified_request_ap_cpu_jtag_debug_module => ap_cpu_data_master_qualified_request_ap_cpu_jtag_debug_module,
      ap_cpu_data_master_qualified_request_clock_crossing_1_s1 => ap_cpu_data_master_qualified_request_clock_crossing_1_s1,
      ap_cpu_data_master_qualified_request_cnApi_Av2Av_0_ap => ap_cpu_data_master_qualified_request_cnApi_Av2Av_0_ap,
      ap_cpu_data_master_qualified_request_jtag_uart_1_avalon_jtag_slave => ap_cpu_data_master_qualified_request_jtag_uart_1_avalon_jtag_slave,
      ap_cpu_data_master_qualified_request_sdram_0_s1 => ap_cpu_data_master_qualified_request_sdram_0_s1,
      ap_cpu_data_master_read => ap_cpu_data_master_read,
      ap_cpu_data_master_read_data_valid_ap_cpu_jtag_debug_module => ap_cpu_data_master_read_data_valid_ap_cpu_jtag_debug_module,
      ap_cpu_data_master_read_data_valid_clock_crossing_1_s1 => ap_cpu_data_master_read_data_valid_clock_crossing_1_s1,
      ap_cpu_data_master_read_data_valid_clock_crossing_1_s1_shift_register => ap_cpu_data_master_read_data_valid_clock_crossing_1_s1_shift_register,
      ap_cpu_data_master_read_data_valid_cnApi_Av2Av_0_ap => ap_cpu_data_master_read_data_valid_cnApi_Av2Av_0_ap,
      ap_cpu_data_master_read_data_valid_jtag_uart_1_avalon_jtag_slave => ap_cpu_data_master_read_data_valid_jtag_uart_1_avalon_jtag_slave,
      ap_cpu_data_master_read_data_valid_sdram_0_s1 => ap_cpu_data_master_read_data_valid_sdram_0_s1,
      ap_cpu_data_master_read_data_valid_sdram_0_s1_shift_register => ap_cpu_data_master_read_data_valid_sdram_0_s1_shift_register,
      ap_cpu_data_master_requests_ap_cpu_jtag_debug_module => ap_cpu_data_master_requests_ap_cpu_jtag_debug_module,
      ap_cpu_data_master_requests_clock_crossing_1_s1 => ap_cpu_data_master_requests_clock_crossing_1_s1,
      ap_cpu_data_master_requests_cnApi_Av2Av_0_ap => ap_cpu_data_master_requests_cnApi_Av2Av_0_ap,
      ap_cpu_data_master_requests_jtag_uart_1_avalon_jtag_slave => ap_cpu_data_master_requests_jtag_uart_1_avalon_jtag_slave,
      ap_cpu_data_master_requests_sdram_0_s1 => ap_cpu_data_master_requests_sdram_0_s1,
      ap_cpu_data_master_write => ap_cpu_data_master_write,
      ap_cpu_jtag_debug_module_readdata_from_sa => ap_cpu_jtag_debug_module_readdata_from_sa,
      clk => internal_clk90Meg,
      clk90Meg => internal_clk90Meg,
      clk90Meg_reset_n => clk90Meg_reset_n,
      clock_crossing_1_s1_readdata_from_sa => clock_crossing_1_s1_readdata_from_sa,
      clock_crossing_1_s1_waitrequest_from_sa => clock_crossing_1_s1_waitrequest_from_sa,
      cnApi_Av2Av_0_ap_readdata_from_sa => cnApi_Av2Av_0_ap_readdata_from_sa,
      cnApi_Av2Av_0_ap_wait_counter_eq_0 => cnApi_Av2Av_0_ap_wait_counter_eq_0,
      d1_ap_cpu_jtag_debug_module_end_xfer => d1_ap_cpu_jtag_debug_module_end_xfer,
      d1_clock_crossing_1_s1_end_xfer => d1_clock_crossing_1_s1_end_xfer,
      d1_cnApi_Av2Av_0_ap_end_xfer => d1_cnApi_Av2Av_0_ap_end_xfer,
      d1_jtag_uart_1_avalon_jtag_slave_end_xfer => d1_jtag_uart_1_avalon_jtag_slave_end_xfer,
      d1_sdram_0_s1_end_xfer => d1_sdram_0_s1_end_xfer,
      jtag_uart_1_avalon_jtag_slave_irq_from_sa => jtag_uart_1_avalon_jtag_slave_irq_from_sa,
      jtag_uart_1_avalon_jtag_slave_readdata_from_sa => jtag_uart_1_avalon_jtag_slave_readdata_from_sa,
      jtag_uart_1_avalon_jtag_slave_waitrequest_from_sa => jtag_uart_1_avalon_jtag_slave_waitrequest_from_sa,
      reset_n => clk90Meg_reset_n,
      sdram_0_s1_readdata_from_sa => sdram_0_s1_readdata_from_sa,
      sdram_0_s1_waitrequest_from_sa => sdram_0_s1_waitrequest_from_sa,
      sync_irq_s1_irq_from_sa => sync_irq_s1_irq_from_sa,
      system_timer_ap_s1_irq_from_sa => system_timer_ap_s1_irq_from_sa
    );


  --the_ap_cpu_instruction_master, which is an e_instance
  the_ap_cpu_instruction_master : ap_cpu_instruction_master_arbitrator
    port map(
      ap_cpu_instruction_master_address_to_slave => ap_cpu_instruction_master_address_to_slave,
      ap_cpu_instruction_master_latency_counter => ap_cpu_instruction_master_latency_counter,
      ap_cpu_instruction_master_readdata => ap_cpu_instruction_master_readdata,
      ap_cpu_instruction_master_readdatavalid => ap_cpu_instruction_master_readdatavalid,
      ap_cpu_instruction_master_waitrequest => ap_cpu_instruction_master_waitrequest,
      ap_cpu_instruction_master_address => ap_cpu_instruction_master_address,
      ap_cpu_instruction_master_granted_ap_cpu_jtag_debug_module => ap_cpu_instruction_master_granted_ap_cpu_jtag_debug_module,
      ap_cpu_instruction_master_granted_sdram_0_s1 => ap_cpu_instruction_master_granted_sdram_0_s1,
      ap_cpu_instruction_master_qualified_request_ap_cpu_jtag_debug_module => ap_cpu_instruction_master_qualified_request_ap_cpu_jtag_debug_module,
      ap_cpu_instruction_master_qualified_request_sdram_0_s1 => ap_cpu_instruction_master_qualified_request_sdram_0_s1,
      ap_cpu_instruction_master_read => ap_cpu_instruction_master_read,
      ap_cpu_instruction_master_read_data_valid_ap_cpu_jtag_debug_module => ap_cpu_instruction_master_read_data_valid_ap_cpu_jtag_debug_module,
      ap_cpu_instruction_master_read_data_valid_sdram_0_s1 => ap_cpu_instruction_master_read_data_valid_sdram_0_s1,
      ap_cpu_instruction_master_read_data_valid_sdram_0_s1_shift_register => ap_cpu_instruction_master_read_data_valid_sdram_0_s1_shift_register,
      ap_cpu_instruction_master_requests_ap_cpu_jtag_debug_module => ap_cpu_instruction_master_requests_ap_cpu_jtag_debug_module,
      ap_cpu_instruction_master_requests_sdram_0_s1 => ap_cpu_instruction_master_requests_sdram_0_s1,
      ap_cpu_jtag_debug_module_readdata_from_sa => ap_cpu_jtag_debug_module_readdata_from_sa,
      clk => internal_clk90Meg,
      d1_ap_cpu_jtag_debug_module_end_xfer => d1_ap_cpu_jtag_debug_module_end_xfer,
      d1_sdram_0_s1_end_xfer => d1_sdram_0_s1_end_xfer,
      reset_n => clk90Meg_reset_n,
      sdram_0_s1_readdata_from_sa => sdram_0_s1_readdata_from_sa,
      sdram_0_s1_waitrequest_from_sa => sdram_0_s1_waitrequest_from_sa
    );


  --the_ap_cpu, which is an e_ptf_instance
  the_ap_cpu : ap_cpu
    port map(
      d_address => ap_cpu_data_master_address,
      d_byteenable => ap_cpu_data_master_byteenable,
      d_read => ap_cpu_data_master_read,
      d_write => ap_cpu_data_master_write,
      d_writedata => ap_cpu_data_master_writedata,
      i_address => ap_cpu_instruction_master_address,
      i_read => ap_cpu_instruction_master_read,
      jtag_debug_module_debugaccess_to_roms => ap_cpu_data_master_debugaccess,
      jtag_debug_module_readdata => ap_cpu_jtag_debug_module_readdata,
      jtag_debug_module_resetrequest => ap_cpu_jtag_debug_module_resetrequest,
      clk => internal_clk90Meg,
      d_irq => ap_cpu_data_master_irq,
      d_readdata => ap_cpu_data_master_readdata,
      d_waitrequest => ap_cpu_data_master_waitrequest,
      i_readdata => ap_cpu_instruction_master_readdata,
      i_readdatavalid => ap_cpu_instruction_master_readdatavalid,
      i_waitrequest => ap_cpu_instruction_master_waitrequest,
      jtag_debug_module_address => ap_cpu_jtag_debug_module_address,
      jtag_debug_module_begintransfer => ap_cpu_jtag_debug_module_begintransfer,
      jtag_debug_module_byteenable => ap_cpu_jtag_debug_module_byteenable,
      jtag_debug_module_debugaccess => ap_cpu_jtag_debug_module_debugaccess,
      jtag_debug_module_select => ap_cpu_jtag_debug_module_chipselect,
      jtag_debug_module_write => ap_cpu_jtag_debug_module_write,
      jtag_debug_module_writedata => ap_cpu_jtag_debug_module_writedata,
      reset_n => ap_cpu_jtag_debug_module_reset_n
    );


  --the_button_pio_s1, which is an e_instance
  the_button_pio_s1 : button_pio_s1_arbitrator
    port map(
      button_pio_s1_address => button_pio_s1_address,
      button_pio_s1_readdata_from_sa => button_pio_s1_readdata_from_sa,
      button_pio_s1_reset_n => button_pio_s1_reset_n,
      clock_crossing_0_m1_granted_button_pio_s1 => clock_crossing_0_m1_granted_button_pio_s1,
      clock_crossing_0_m1_qualified_request_button_pio_s1 => clock_crossing_0_m1_qualified_request_button_pio_s1,
      clock_crossing_0_m1_read_data_valid_button_pio_s1 => clock_crossing_0_m1_read_data_valid_button_pio_s1,
      clock_crossing_0_m1_requests_button_pio_s1 => clock_crossing_0_m1_requests_button_pio_s1,
      d1_button_pio_s1_end_xfer => d1_button_pio_s1_end_xfer,
      button_pio_s1_readdata => button_pio_s1_readdata,
      clk => internal_clk50Meg,
      clock_crossing_0_m1_address_to_slave => clock_crossing_0_m1_address_to_slave,
      clock_crossing_0_m1_latency_counter => clock_crossing_0_m1_latency_counter,
      clock_crossing_0_m1_nativeaddress => clock_crossing_0_m1_nativeaddress,
      clock_crossing_0_m1_read => clock_crossing_0_m1_read,
      clock_crossing_0_m1_write => clock_crossing_0_m1_write,
      reset_n => clk50Meg_reset_n
    );


  --the_button_pio, which is an e_ptf_instance
  the_button_pio : button_pio
    port map(
      readdata => button_pio_s1_readdata,
      address => button_pio_s1_address,
      clk => internal_clk50Meg,
      in_port => in_port_to_the_button_pio,
      reset_n => button_pio_s1_reset_n
    );


  --the_clock_crossing_0_s1, which is an e_instance
  the_clock_crossing_0_s1 : clock_crossing_0_s1_arbitrator
    port map(
      clock_crossing_0_s1_address => clock_crossing_0_s1_address,
      clock_crossing_0_s1_byteenable => clock_crossing_0_s1_byteenable,
      clock_crossing_0_s1_endofpacket_from_sa => clock_crossing_0_s1_endofpacket_from_sa,
      clock_crossing_0_s1_nativeaddress => clock_crossing_0_s1_nativeaddress,
      clock_crossing_0_s1_read => clock_crossing_0_s1_read,
      clock_crossing_0_s1_readdata_from_sa => clock_crossing_0_s1_readdata_from_sa,
      clock_crossing_0_s1_reset_n => clock_crossing_0_s1_reset_n,
      clock_crossing_0_s1_waitrequest_from_sa => clock_crossing_0_s1_waitrequest_from_sa,
      clock_crossing_0_s1_write => clock_crossing_0_s1_write,
      clock_crossing_0_s1_writedata => clock_crossing_0_s1_writedata,
      d1_clock_crossing_0_s1_end_xfer => d1_clock_crossing_0_s1_end_xfer,
      pcp_cpu_data_master_granted_clock_crossing_0_s1 => pcp_cpu_data_master_granted_clock_crossing_0_s1,
      pcp_cpu_data_master_qualified_request_clock_crossing_0_s1 => pcp_cpu_data_master_qualified_request_clock_crossing_0_s1,
      pcp_cpu_data_master_read_data_valid_clock_crossing_0_s1 => pcp_cpu_data_master_read_data_valid_clock_crossing_0_s1,
      pcp_cpu_data_master_read_data_valid_clock_crossing_0_s1_shift_register => pcp_cpu_data_master_read_data_valid_clock_crossing_0_s1_shift_register,
      pcp_cpu_data_master_requests_clock_crossing_0_s1 => pcp_cpu_data_master_requests_clock_crossing_0_s1,
      clk => internal_clk90Meg,
      clock_crossing_0_s1_endofpacket => clock_crossing_0_s1_endofpacket,
      clock_crossing_0_s1_readdata => clock_crossing_0_s1_readdata,
      clock_crossing_0_s1_readdatavalid => clock_crossing_0_s1_readdatavalid,
      clock_crossing_0_s1_waitrequest => clock_crossing_0_s1_waitrequest,
      pcp_cpu_data_master_address_to_slave => pcp_cpu_data_master_address_to_slave,
      pcp_cpu_data_master_byteenable => pcp_cpu_data_master_byteenable,
      pcp_cpu_data_master_read => pcp_cpu_data_master_read,
      pcp_cpu_data_master_waitrequest => pcp_cpu_data_master_waitrequest,
      pcp_cpu_data_master_write => pcp_cpu_data_master_write,
      pcp_cpu_data_master_writedata => pcp_cpu_data_master_writedata,
      reset_n => clk90Meg_reset_n
    );


  --the_clock_crossing_0_m1, which is an e_instance
  the_clock_crossing_0_m1 : clock_crossing_0_m1_arbitrator
    port map(
      clock_crossing_0_m1_address_to_slave => clock_crossing_0_m1_address_to_slave,
      clock_crossing_0_m1_latency_counter => clock_crossing_0_m1_latency_counter,
      clock_crossing_0_m1_readdata => clock_crossing_0_m1_readdata,
      clock_crossing_0_m1_readdatavalid => clock_crossing_0_m1_readdatavalid,
      clock_crossing_0_m1_reset_n => clock_crossing_0_m1_reset_n,
      clock_crossing_0_m1_waitrequest => clock_crossing_0_m1_waitrequest,
      button_pio_s1_readdata_from_sa => button_pio_s1_readdata_from_sa,
      clk => internal_clk50Meg,
      clock_crossing_0_m1_address => clock_crossing_0_m1_address,
      clock_crossing_0_m1_byteenable => clock_crossing_0_m1_byteenable,
      clock_crossing_0_m1_granted_button_pio_s1 => clock_crossing_0_m1_granted_button_pio_s1,
      clock_crossing_0_m1_granted_irq_gen_s1 => clock_crossing_0_m1_granted_irq_gen_s1,
      clock_crossing_0_m1_granted_status_led_pio_s1 => clock_crossing_0_m1_granted_status_led_pio_s1,
      clock_crossing_0_m1_granted_sysid_control_slave => clock_crossing_0_m1_granted_sysid_control_slave,
      clock_crossing_0_m1_granted_system_timer_s1 => clock_crossing_0_m1_granted_system_timer_s1,
      clock_crossing_0_m1_qualified_request_button_pio_s1 => clock_crossing_0_m1_qualified_request_button_pio_s1,
      clock_crossing_0_m1_qualified_request_irq_gen_s1 => clock_crossing_0_m1_qualified_request_irq_gen_s1,
      clock_crossing_0_m1_qualified_request_status_led_pio_s1 => clock_crossing_0_m1_qualified_request_status_led_pio_s1,
      clock_crossing_0_m1_qualified_request_sysid_control_slave => clock_crossing_0_m1_qualified_request_sysid_control_slave,
      clock_crossing_0_m1_qualified_request_system_timer_s1 => clock_crossing_0_m1_qualified_request_system_timer_s1,
      clock_crossing_0_m1_read => clock_crossing_0_m1_read,
      clock_crossing_0_m1_read_data_valid_button_pio_s1 => clock_crossing_0_m1_read_data_valid_button_pio_s1,
      clock_crossing_0_m1_read_data_valid_irq_gen_s1 => clock_crossing_0_m1_read_data_valid_irq_gen_s1,
      clock_crossing_0_m1_read_data_valid_status_led_pio_s1 => clock_crossing_0_m1_read_data_valid_status_led_pio_s1,
      clock_crossing_0_m1_read_data_valid_sysid_control_slave => clock_crossing_0_m1_read_data_valid_sysid_control_slave,
      clock_crossing_0_m1_read_data_valid_system_timer_s1 => clock_crossing_0_m1_read_data_valid_system_timer_s1,
      clock_crossing_0_m1_requests_button_pio_s1 => clock_crossing_0_m1_requests_button_pio_s1,
      clock_crossing_0_m1_requests_irq_gen_s1 => clock_crossing_0_m1_requests_irq_gen_s1,
      clock_crossing_0_m1_requests_status_led_pio_s1 => clock_crossing_0_m1_requests_status_led_pio_s1,
      clock_crossing_0_m1_requests_sysid_control_slave => clock_crossing_0_m1_requests_sysid_control_slave,
      clock_crossing_0_m1_requests_system_timer_s1 => clock_crossing_0_m1_requests_system_timer_s1,
      clock_crossing_0_m1_write => clock_crossing_0_m1_write,
      clock_crossing_0_m1_writedata => clock_crossing_0_m1_writedata,
      d1_button_pio_s1_end_xfer => d1_button_pio_s1_end_xfer,
      d1_irq_gen_s1_end_xfer => d1_irq_gen_s1_end_xfer,
      d1_status_led_pio_s1_end_xfer => d1_status_led_pio_s1_end_xfer,
      d1_sysid_control_slave_end_xfer => d1_sysid_control_slave_end_xfer,
      d1_system_timer_s1_end_xfer => d1_system_timer_s1_end_xfer,
      irq_gen_s1_readdata_from_sa => irq_gen_s1_readdata_from_sa,
      reset_n => clk50Meg_reset_n,
      status_led_pio_s1_readdata_from_sa => status_led_pio_s1_readdata_from_sa,
      sysid_control_slave_readdata_from_sa => sysid_control_slave_readdata_from_sa,
      system_timer_s1_readdata_from_sa => system_timer_s1_readdata_from_sa
    );


  --the_clock_crossing_0, which is an e_ptf_instance
  the_clock_crossing_0 : clock_crossing_0
    port map(
      master_address => clock_crossing_0_m1_address,
      master_byteenable => clock_crossing_0_m1_byteenable,
      master_nativeaddress => clock_crossing_0_m1_nativeaddress,
      master_read => clock_crossing_0_m1_read,
      master_write => clock_crossing_0_m1_write,
      master_writedata => clock_crossing_0_m1_writedata,
      slave_endofpacket => clock_crossing_0_s1_endofpacket,
      slave_readdata => clock_crossing_0_s1_readdata,
      slave_readdatavalid => clock_crossing_0_s1_readdatavalid,
      slave_waitrequest => clock_crossing_0_s1_waitrequest,
      master_clk => internal_clk50Meg,
      master_endofpacket => clock_crossing_0_m1_endofpacket,
      master_readdata => clock_crossing_0_m1_readdata,
      master_readdatavalid => clock_crossing_0_m1_readdatavalid,
      master_reset_n => clock_crossing_0_m1_reset_n,
      master_waitrequest => clock_crossing_0_m1_waitrequest,
      slave_address => clock_crossing_0_s1_address,
      slave_byteenable => clock_crossing_0_s1_byteenable,
      slave_clk => internal_clk90Meg,
      slave_nativeaddress => clock_crossing_0_s1_nativeaddress,
      slave_read => clock_crossing_0_s1_read,
      slave_reset_n => clock_crossing_0_s1_reset_n,
      slave_write => clock_crossing_0_s1_write,
      slave_writedata => clock_crossing_0_s1_writedata
    );


  --the_clock_crossing_1_s1, which is an e_instance
  the_clock_crossing_1_s1 : clock_crossing_1_s1_arbitrator
    port map(
      ap_cpu_data_master_granted_clock_crossing_1_s1 => ap_cpu_data_master_granted_clock_crossing_1_s1,
      ap_cpu_data_master_qualified_request_clock_crossing_1_s1 => ap_cpu_data_master_qualified_request_clock_crossing_1_s1,
      ap_cpu_data_master_read_data_valid_clock_crossing_1_s1 => ap_cpu_data_master_read_data_valid_clock_crossing_1_s1,
      ap_cpu_data_master_read_data_valid_clock_crossing_1_s1_shift_register => ap_cpu_data_master_read_data_valid_clock_crossing_1_s1_shift_register,
      ap_cpu_data_master_requests_clock_crossing_1_s1 => ap_cpu_data_master_requests_clock_crossing_1_s1,
      clock_crossing_1_s1_address => clock_crossing_1_s1_address,
      clock_crossing_1_s1_byteenable => clock_crossing_1_s1_byteenable,
      clock_crossing_1_s1_endofpacket_from_sa => clock_crossing_1_s1_endofpacket_from_sa,
      clock_crossing_1_s1_nativeaddress => clock_crossing_1_s1_nativeaddress,
      clock_crossing_1_s1_read => clock_crossing_1_s1_read,
      clock_crossing_1_s1_readdata_from_sa => clock_crossing_1_s1_readdata_from_sa,
      clock_crossing_1_s1_reset_n => clock_crossing_1_s1_reset_n,
      clock_crossing_1_s1_waitrequest_from_sa => clock_crossing_1_s1_waitrequest_from_sa,
      clock_crossing_1_s1_write => clock_crossing_1_s1_write,
      clock_crossing_1_s1_writedata => clock_crossing_1_s1_writedata,
      d1_clock_crossing_1_s1_end_xfer => d1_clock_crossing_1_s1_end_xfer,
      ap_cpu_data_master_address_to_slave => ap_cpu_data_master_address_to_slave,
      ap_cpu_data_master_byteenable => ap_cpu_data_master_byteenable,
      ap_cpu_data_master_read => ap_cpu_data_master_read,
      ap_cpu_data_master_waitrequest => ap_cpu_data_master_waitrequest,
      ap_cpu_data_master_write => ap_cpu_data_master_write,
      ap_cpu_data_master_writedata => ap_cpu_data_master_writedata,
      clk => internal_clk90Meg,
      clock_crossing_1_s1_endofpacket => clock_crossing_1_s1_endofpacket,
      clock_crossing_1_s1_readdata => clock_crossing_1_s1_readdata,
      clock_crossing_1_s1_readdatavalid => clock_crossing_1_s1_readdatavalid,
      clock_crossing_1_s1_waitrequest => clock_crossing_1_s1_waitrequest,
      reset_n => clk90Meg_reset_n
    );


  --the_clock_crossing_1_m1, which is an e_instance
  the_clock_crossing_1_m1 : clock_crossing_1_m1_arbitrator
    port map(
      clock_crossing_1_m1_address_to_slave => clock_crossing_1_m1_address_to_slave,
      clock_crossing_1_m1_latency_counter => clock_crossing_1_m1_latency_counter,
      clock_crossing_1_m1_readdata => clock_crossing_1_m1_readdata,
      clock_crossing_1_m1_readdatavalid => clock_crossing_1_m1_readdatavalid,
      clock_crossing_1_m1_reset_n => clock_crossing_1_m1_reset_n,
      clock_crossing_1_m1_waitrequest => clock_crossing_1_m1_waitrequest,
      clk => internal_clk50Meg,
      clock_crossing_1_m1_address => clock_crossing_1_m1_address,
      clock_crossing_1_m1_byteenable => clock_crossing_1_m1_byteenable,
      clock_crossing_1_m1_granted_digio_pio_s1 => clock_crossing_1_m1_granted_digio_pio_s1,
      clock_crossing_1_m1_granted_node_switch_pio_s1 => clock_crossing_1_m1_granted_node_switch_pio_s1,
      clock_crossing_1_m1_granted_portconf_pio_s1 => clock_crossing_1_m1_granted_portconf_pio_s1,
      clock_crossing_1_m1_granted_sync_irq_s1 => clock_crossing_1_m1_granted_sync_irq_s1,
      clock_crossing_1_m1_granted_sysid_control_slave => clock_crossing_1_m1_granted_sysid_control_slave,
      clock_crossing_1_m1_granted_system_timer_ap_s1 => clock_crossing_1_m1_granted_system_timer_ap_s1,
      clock_crossing_1_m1_qualified_request_digio_pio_s1 => clock_crossing_1_m1_qualified_request_digio_pio_s1,
      clock_crossing_1_m1_qualified_request_node_switch_pio_s1 => clock_crossing_1_m1_qualified_request_node_switch_pio_s1,
      clock_crossing_1_m1_qualified_request_portconf_pio_s1 => clock_crossing_1_m1_qualified_request_portconf_pio_s1,
      clock_crossing_1_m1_qualified_request_sync_irq_s1 => clock_crossing_1_m1_qualified_request_sync_irq_s1,
      clock_crossing_1_m1_qualified_request_sysid_control_slave => clock_crossing_1_m1_qualified_request_sysid_control_slave,
      clock_crossing_1_m1_qualified_request_system_timer_ap_s1 => clock_crossing_1_m1_qualified_request_system_timer_ap_s1,
      clock_crossing_1_m1_read => clock_crossing_1_m1_read,
      clock_crossing_1_m1_read_data_valid_digio_pio_s1 => clock_crossing_1_m1_read_data_valid_digio_pio_s1,
      clock_crossing_1_m1_read_data_valid_node_switch_pio_s1 => clock_crossing_1_m1_read_data_valid_node_switch_pio_s1,
      clock_crossing_1_m1_read_data_valid_portconf_pio_s1 => clock_crossing_1_m1_read_data_valid_portconf_pio_s1,
      clock_crossing_1_m1_read_data_valid_sync_irq_s1 => clock_crossing_1_m1_read_data_valid_sync_irq_s1,
      clock_crossing_1_m1_read_data_valid_sysid_control_slave => clock_crossing_1_m1_read_data_valid_sysid_control_slave,
      clock_crossing_1_m1_read_data_valid_system_timer_ap_s1 => clock_crossing_1_m1_read_data_valid_system_timer_ap_s1,
      clock_crossing_1_m1_requests_digio_pio_s1 => clock_crossing_1_m1_requests_digio_pio_s1,
      clock_crossing_1_m1_requests_node_switch_pio_s1 => clock_crossing_1_m1_requests_node_switch_pio_s1,
      clock_crossing_1_m1_requests_portconf_pio_s1 => clock_crossing_1_m1_requests_portconf_pio_s1,
      clock_crossing_1_m1_requests_sync_irq_s1 => clock_crossing_1_m1_requests_sync_irq_s1,
      clock_crossing_1_m1_requests_sysid_control_slave => clock_crossing_1_m1_requests_sysid_control_slave,
      clock_crossing_1_m1_requests_system_timer_ap_s1 => clock_crossing_1_m1_requests_system_timer_ap_s1,
      clock_crossing_1_m1_write => clock_crossing_1_m1_write,
      clock_crossing_1_m1_writedata => clock_crossing_1_m1_writedata,
      d1_digio_pio_s1_end_xfer => d1_digio_pio_s1_end_xfer,
      d1_node_switch_pio_s1_end_xfer => d1_node_switch_pio_s1_end_xfer,
      d1_portconf_pio_s1_end_xfer => d1_portconf_pio_s1_end_xfer,
      d1_sync_irq_s1_end_xfer => d1_sync_irq_s1_end_xfer,
      d1_sysid_control_slave_end_xfer => d1_sysid_control_slave_end_xfer,
      d1_system_timer_ap_s1_end_xfer => d1_system_timer_ap_s1_end_xfer,
      digio_pio_s1_readdata_from_sa => digio_pio_s1_readdata_from_sa,
      node_switch_pio_s1_readdata_from_sa => node_switch_pio_s1_readdata_from_sa,
      portconf_pio_s1_readdata_from_sa => portconf_pio_s1_readdata_from_sa,
      reset_n => clk50Meg_reset_n,
      sync_irq_s1_readdata_from_sa => sync_irq_s1_readdata_from_sa,
      sysid_control_slave_readdata_from_sa => sysid_control_slave_readdata_from_sa,
      system_timer_ap_s1_readdata_from_sa => system_timer_ap_s1_readdata_from_sa
    );


  --the_clock_crossing_1, which is an e_ptf_instance
  the_clock_crossing_1 : clock_crossing_1
    port map(
      master_address => clock_crossing_1_m1_address,
      master_byteenable => clock_crossing_1_m1_byteenable,
      master_nativeaddress => clock_crossing_1_m1_nativeaddress,
      master_read => clock_crossing_1_m1_read,
      master_write => clock_crossing_1_m1_write,
      master_writedata => clock_crossing_1_m1_writedata,
      slave_endofpacket => clock_crossing_1_s1_endofpacket,
      slave_readdata => clock_crossing_1_s1_readdata,
      slave_readdatavalid => clock_crossing_1_s1_readdatavalid,
      slave_waitrequest => clock_crossing_1_s1_waitrequest,
      master_clk => internal_clk50Meg,
      master_endofpacket => clock_crossing_1_m1_endofpacket,
      master_readdata => clock_crossing_1_m1_readdata,
      master_readdatavalid => clock_crossing_1_m1_readdatavalid,
      master_reset_n => clock_crossing_1_m1_reset_n,
      master_waitrequest => clock_crossing_1_m1_waitrequest,
      slave_address => clock_crossing_1_s1_address,
      slave_byteenable => clock_crossing_1_s1_byteenable,
      slave_clk => internal_clk90Meg,
      slave_nativeaddress => clock_crossing_1_s1_nativeaddress,
      slave_read => clock_crossing_1_s1_read,
      slave_reset_n => clock_crossing_1_s1_reset_n,
      slave_write => clock_crossing_1_s1_write,
      slave_writedata => clock_crossing_1_s1_writedata
    );


  --the_cnApi_Av2Av_0_ap, which is an e_instance
  the_cnApi_Av2Av_0_ap : cnApi_Av2Av_0_ap_arbitrator
    port map(
      ap_cpu_data_master_granted_cnApi_Av2Av_0_ap => ap_cpu_data_master_granted_cnApi_Av2Av_0_ap,
      ap_cpu_data_master_qualified_request_cnApi_Av2Av_0_ap => ap_cpu_data_master_qualified_request_cnApi_Av2Av_0_ap,
      ap_cpu_data_master_read_data_valid_cnApi_Av2Av_0_ap => ap_cpu_data_master_read_data_valid_cnApi_Av2Av_0_ap,
      ap_cpu_data_master_requests_cnApi_Av2Av_0_ap => ap_cpu_data_master_requests_cnApi_Av2Av_0_ap,
      cnApi_Av2Av_0_ap_address => cnApi_Av2Av_0_ap_address,
      cnApi_Av2Av_0_ap_byteenable => cnApi_Av2Av_0_ap_byteenable,
      cnApi_Av2Av_0_ap_chipselect => cnApi_Av2Av_0_ap_chipselect,
      cnApi_Av2Av_0_ap_read => cnApi_Av2Av_0_ap_read,
      cnApi_Av2Av_0_ap_readdata_from_sa => cnApi_Av2Av_0_ap_readdata_from_sa,
      cnApi_Av2Av_0_ap_reset => cnApi_Av2Av_0_ap_reset,
      cnApi_Av2Av_0_ap_wait_counter_eq_0 => cnApi_Av2Av_0_ap_wait_counter_eq_0,
      cnApi_Av2Av_0_ap_write => cnApi_Av2Av_0_ap_write,
      cnApi_Av2Av_0_ap_writedata => cnApi_Av2Av_0_ap_writedata,
      d1_cnApi_Av2Av_0_ap_end_xfer => d1_cnApi_Av2Av_0_ap_end_xfer,
      ap_cpu_data_master_address_to_slave => ap_cpu_data_master_address_to_slave,
      ap_cpu_data_master_byteenable => ap_cpu_data_master_byteenable,
      ap_cpu_data_master_read => ap_cpu_data_master_read,
      ap_cpu_data_master_waitrequest => ap_cpu_data_master_waitrequest,
      ap_cpu_data_master_write => ap_cpu_data_master_write,
      ap_cpu_data_master_writedata => ap_cpu_data_master_writedata,
      clk => internal_clk90Meg,
      cnApi_Av2Av_0_ap_readdata => cnApi_Av2Av_0_ap_readdata,
      reset_n => clk90Meg_reset_n
    );


  --the_cnApi_Av2Av_0_pcp, which is an e_instance
  the_cnApi_Av2Av_0_pcp : cnApi_Av2Av_0_pcp_arbitrator
    port map(
      cnApi_Av2Av_0_pcp_address => cnApi_Av2Av_0_pcp_address,
      cnApi_Av2Av_0_pcp_byteenable => cnApi_Av2Av_0_pcp_byteenable,
      cnApi_Av2Av_0_pcp_chipselect => cnApi_Av2Av_0_pcp_chipselect,
      cnApi_Av2Av_0_pcp_read => cnApi_Av2Av_0_pcp_read,
      cnApi_Av2Av_0_pcp_readdata_from_sa => cnApi_Av2Av_0_pcp_readdata_from_sa,
      cnApi_Av2Av_0_pcp_reset => cnApi_Av2Av_0_pcp_reset,
      cnApi_Av2Av_0_pcp_wait_counter_eq_0 => cnApi_Av2Av_0_pcp_wait_counter_eq_0,
      cnApi_Av2Av_0_pcp_write => cnApi_Av2Av_0_pcp_write,
      cnApi_Av2Av_0_pcp_writedata => cnApi_Av2Av_0_pcp_writedata,
      d1_cnApi_Av2Av_0_pcp_end_xfer => d1_cnApi_Av2Av_0_pcp_end_xfer,
      pcp_cpu_data_master_granted_cnApi_Av2Av_0_pcp => pcp_cpu_data_master_granted_cnApi_Av2Av_0_pcp,
      pcp_cpu_data_master_qualified_request_cnApi_Av2Av_0_pcp => pcp_cpu_data_master_qualified_request_cnApi_Av2Av_0_pcp,
      pcp_cpu_data_master_read_data_valid_cnApi_Av2Av_0_pcp => pcp_cpu_data_master_read_data_valid_cnApi_Av2Av_0_pcp,
      pcp_cpu_data_master_requests_cnApi_Av2Av_0_pcp => pcp_cpu_data_master_requests_cnApi_Av2Av_0_pcp,
      clk => internal_clk90Meg,
      cnApi_Av2Av_0_pcp_readdata => cnApi_Av2Av_0_pcp_readdata,
      pcp_cpu_data_master_address_to_slave => pcp_cpu_data_master_address_to_slave,
      pcp_cpu_data_master_byteenable => pcp_cpu_data_master_byteenable,
      pcp_cpu_data_master_read => pcp_cpu_data_master_read,
      pcp_cpu_data_master_waitrequest => pcp_cpu_data_master_waitrequest,
      pcp_cpu_data_master_write => pcp_cpu_data_master_write,
      pcp_cpu_data_master_writedata => pcp_cpu_data_master_writedata,
      reset_n => clk90Meg_reset_n
    );


  --the_cnApi_Av2Av_0, which is an e_ptf_instance
  the_cnApi_Av2Av_0 : cnApi_Av2Av_0
    port map(
      ap_readdata => cnApi_Av2Av_0_ap_readdata,
      pcp_readdata => cnApi_Av2Av_0_pcp_readdata,
      ap_Clk => internal_clk90Meg,
      ap_Reset => cnApi_Av2Av_0_ap_reset,
      ap_address => cnApi_Av2Av_0_ap_address,
      ap_byteenable => cnApi_Av2Av_0_ap_byteenable,
      ap_chipselect => cnApi_Av2Av_0_ap_chipselect,
      ap_read => cnApi_Av2Av_0_ap_read,
      ap_write => cnApi_Av2Av_0_ap_write,
      ap_writedata => cnApi_Av2Av_0_ap_writedata,
      pcp_Clk => internal_clk90Meg,
      pcp_Reset => cnApi_Av2Av_0_pcp_reset,
      pcp_address => cnApi_Av2Av_0_pcp_address,
      pcp_byteenable => cnApi_Av2Av_0_pcp_byteenable,
      pcp_chipselect => cnApi_Av2Av_0_pcp_chipselect,
      pcp_read => cnApi_Av2Av_0_pcp_read,
      pcp_write => cnApi_Av2Av_0_pcp_write,
      pcp_writedata => cnApi_Av2Av_0_pcp_writedata
    );


  --the_digio_pio_s1, which is an e_instance
  the_digio_pio_s1 : digio_pio_s1_arbitrator
    port map(
      clock_crossing_1_m1_granted_digio_pio_s1 => clock_crossing_1_m1_granted_digio_pio_s1,
      clock_crossing_1_m1_qualified_request_digio_pio_s1 => clock_crossing_1_m1_qualified_request_digio_pio_s1,
      clock_crossing_1_m1_read_data_valid_digio_pio_s1 => clock_crossing_1_m1_read_data_valid_digio_pio_s1,
      clock_crossing_1_m1_requests_digio_pio_s1 => clock_crossing_1_m1_requests_digio_pio_s1,
      d1_digio_pio_s1_end_xfer => d1_digio_pio_s1_end_xfer,
      digio_pio_s1_address => digio_pio_s1_address,
      digio_pio_s1_chipselect => digio_pio_s1_chipselect,
      digio_pio_s1_readdata_from_sa => digio_pio_s1_readdata_from_sa,
      digio_pio_s1_reset_n => digio_pio_s1_reset_n,
      digio_pio_s1_write_n => digio_pio_s1_write_n,
      digio_pio_s1_writedata => digio_pio_s1_writedata,
      clk => internal_clk50Meg,
      clock_crossing_1_m1_address_to_slave => clock_crossing_1_m1_address_to_slave,
      clock_crossing_1_m1_latency_counter => clock_crossing_1_m1_latency_counter,
      clock_crossing_1_m1_nativeaddress => clock_crossing_1_m1_nativeaddress,
      clock_crossing_1_m1_read => clock_crossing_1_m1_read,
      clock_crossing_1_m1_write => clock_crossing_1_m1_write,
      clock_crossing_1_m1_writedata => clock_crossing_1_m1_writedata,
      digio_pio_s1_readdata => digio_pio_s1_readdata,
      reset_n => clk50Meg_reset_n
    );


  --the_digio_pio, which is an e_ptf_instance
  the_digio_pio : digio_pio
    port map(
      bidir_port => bidir_port_to_and_from_the_digio_pio,
      readdata => digio_pio_s1_readdata,
      address => digio_pio_s1_address,
      chipselect => digio_pio_s1_chipselect,
      clk => internal_clk50Meg,
      reset_n => digio_pio_s1_reset_n,
      write_n => digio_pio_s1_write_n,
      writedata => digio_pio_s1_writedata
    );


  --the_epcs_flash_controller_0_epcs_control_port, which is an e_instance
  the_epcs_flash_controller_0_epcs_control_port : epcs_flash_controller_0_epcs_control_port_arbitrator
    port map(
      d1_epcs_flash_controller_0_epcs_control_port_end_xfer => d1_epcs_flash_controller_0_epcs_control_port_end_xfer,
      epcs_flash_controller_0_epcs_control_port_address => epcs_flash_controller_0_epcs_control_port_address,
      epcs_flash_controller_0_epcs_control_port_chipselect => epcs_flash_controller_0_epcs_control_port_chipselect,
      epcs_flash_controller_0_epcs_control_port_dataavailable_from_sa => epcs_flash_controller_0_epcs_control_port_dataavailable_from_sa,
      epcs_flash_controller_0_epcs_control_port_endofpacket_from_sa => epcs_flash_controller_0_epcs_control_port_endofpacket_from_sa,
      epcs_flash_controller_0_epcs_control_port_irq_from_sa => epcs_flash_controller_0_epcs_control_port_irq_from_sa,
      epcs_flash_controller_0_epcs_control_port_read_n => epcs_flash_controller_0_epcs_control_port_read_n,
      epcs_flash_controller_0_epcs_control_port_readdata_from_sa => epcs_flash_controller_0_epcs_control_port_readdata_from_sa,
      epcs_flash_controller_0_epcs_control_port_readyfordata_from_sa => epcs_flash_controller_0_epcs_control_port_readyfordata_from_sa,
      epcs_flash_controller_0_epcs_control_port_reset_n => epcs_flash_controller_0_epcs_control_port_reset_n,
      epcs_flash_controller_0_epcs_control_port_write_n => epcs_flash_controller_0_epcs_control_port_write_n,
      epcs_flash_controller_0_epcs_control_port_writedata => epcs_flash_controller_0_epcs_control_port_writedata,
      pcp_cpu_data_master_granted_epcs_flash_controller_0_epcs_control_port => pcp_cpu_data_master_granted_epcs_flash_controller_0_epcs_control_port,
      pcp_cpu_data_master_qualified_request_epcs_flash_controller_0_epcs_control_port => pcp_cpu_data_master_qualified_request_epcs_flash_controller_0_epcs_control_port,
      pcp_cpu_data_master_read_data_valid_epcs_flash_controller_0_epcs_control_port => pcp_cpu_data_master_read_data_valid_epcs_flash_controller_0_epcs_control_port,
      pcp_cpu_data_master_requests_epcs_flash_controller_0_epcs_control_port => pcp_cpu_data_master_requests_epcs_flash_controller_0_epcs_control_port,
      pcp_cpu_instruction_master_granted_epcs_flash_controller_0_epcs_control_port => pcp_cpu_instruction_master_granted_epcs_flash_controller_0_epcs_control_port,
      pcp_cpu_instruction_master_qualified_request_epcs_flash_controller_0_epcs_control_port => pcp_cpu_instruction_master_qualified_request_epcs_flash_controller_0_epcs_control_port,
      pcp_cpu_instruction_master_read_data_valid_epcs_flash_controller_0_epcs_control_port => pcp_cpu_instruction_master_read_data_valid_epcs_flash_controller_0_epcs_control_port,
      pcp_cpu_instruction_master_requests_epcs_flash_controller_0_epcs_control_port => pcp_cpu_instruction_master_requests_epcs_flash_controller_0_epcs_control_port,
      clk => internal_clk90Meg,
      epcs_flash_controller_0_epcs_control_port_dataavailable => epcs_flash_controller_0_epcs_control_port_dataavailable,
      epcs_flash_controller_0_epcs_control_port_endofpacket => epcs_flash_controller_0_epcs_control_port_endofpacket,
      epcs_flash_controller_0_epcs_control_port_irq => epcs_flash_controller_0_epcs_control_port_irq,
      epcs_flash_controller_0_epcs_control_port_readdata => epcs_flash_controller_0_epcs_control_port_readdata,
      epcs_flash_controller_0_epcs_control_port_readyfordata => epcs_flash_controller_0_epcs_control_port_readyfordata,
      pcp_cpu_data_master_address_to_slave => pcp_cpu_data_master_address_to_slave,
      pcp_cpu_data_master_read => pcp_cpu_data_master_read,
      pcp_cpu_data_master_write => pcp_cpu_data_master_write,
      pcp_cpu_data_master_writedata => pcp_cpu_data_master_writedata,
      pcp_cpu_instruction_master_address_to_slave => pcp_cpu_instruction_master_address_to_slave,
      pcp_cpu_instruction_master_latency_counter => pcp_cpu_instruction_master_latency_counter,
      pcp_cpu_instruction_master_read => pcp_cpu_instruction_master_read,
      reset_n => clk90Meg_reset_n
    );


  --the_epcs_flash_controller_0, which is an e_ptf_instance
  the_epcs_flash_controller_0 : epcs_flash_controller_0
    port map(
      dataavailable => epcs_flash_controller_0_epcs_control_port_dataavailable,
      dclk => internal_dclk_from_the_epcs_flash_controller_0,
      endofpacket => epcs_flash_controller_0_epcs_control_port_endofpacket,
      irq => epcs_flash_controller_0_epcs_control_port_irq,
      readdata => epcs_flash_controller_0_epcs_control_port_readdata,
      readyfordata => epcs_flash_controller_0_epcs_control_port_readyfordata,
      sce => internal_sce_from_the_epcs_flash_controller_0,
      sdo => internal_sdo_from_the_epcs_flash_controller_0,
      address => epcs_flash_controller_0_epcs_control_port_address,
      chipselect => epcs_flash_controller_0_epcs_control_port_chipselect,
      clk => internal_clk90Meg,
      data0 => data0_to_the_epcs_flash_controller_0,
      read_n => epcs_flash_controller_0_epcs_control_port_read_n,
      reset_n => epcs_flash_controller_0_epcs_control_port_reset_n,
      write_n => epcs_flash_controller_0_epcs_control_port_write_n,
      writedata => epcs_flash_controller_0_epcs_control_port_writedata
    );


  --the_irq_gen_s1, which is an e_instance
  the_irq_gen_s1 : irq_gen_s1_arbitrator
    port map(
      clock_crossing_0_m1_granted_irq_gen_s1 => clock_crossing_0_m1_granted_irq_gen_s1,
      clock_crossing_0_m1_qualified_request_irq_gen_s1 => clock_crossing_0_m1_qualified_request_irq_gen_s1,
      clock_crossing_0_m1_read_data_valid_irq_gen_s1 => clock_crossing_0_m1_read_data_valid_irq_gen_s1,
      clock_crossing_0_m1_requests_irq_gen_s1 => clock_crossing_0_m1_requests_irq_gen_s1,
      d1_irq_gen_s1_end_xfer => d1_irq_gen_s1_end_xfer,
      irq_gen_s1_address => irq_gen_s1_address,
      irq_gen_s1_chipselect => irq_gen_s1_chipselect,
      irq_gen_s1_readdata_from_sa => irq_gen_s1_readdata_from_sa,
      irq_gen_s1_reset_n => irq_gen_s1_reset_n,
      irq_gen_s1_write_n => irq_gen_s1_write_n,
      irq_gen_s1_writedata => irq_gen_s1_writedata,
      clk => internal_clk50Meg,
      clock_crossing_0_m1_address_to_slave => clock_crossing_0_m1_address_to_slave,
      clock_crossing_0_m1_latency_counter => clock_crossing_0_m1_latency_counter,
      clock_crossing_0_m1_nativeaddress => clock_crossing_0_m1_nativeaddress,
      clock_crossing_0_m1_read => clock_crossing_0_m1_read,
      clock_crossing_0_m1_write => clock_crossing_0_m1_write,
      clock_crossing_0_m1_writedata => clock_crossing_0_m1_writedata,
      irq_gen_s1_readdata => irq_gen_s1_readdata,
      reset_n => clk50Meg_reset_n
    );


  --the_irq_gen, which is an e_ptf_instance
  the_irq_gen : irq_gen
    port map(
      out_port => internal_out_port_from_the_irq_gen,
      readdata => irq_gen_s1_readdata,
      address => irq_gen_s1_address,
      chipselect => irq_gen_s1_chipselect,
      clk => internal_clk50Meg,
      reset_n => irq_gen_s1_reset_n,
      write_n => irq_gen_s1_write_n,
      writedata => irq_gen_s1_writedata
    );


  --the_jtag_uart_0_avalon_jtag_slave, which is an e_instance
  the_jtag_uart_0_avalon_jtag_slave : jtag_uart_0_avalon_jtag_slave_arbitrator
    port map(
      d1_jtag_uart_0_avalon_jtag_slave_end_xfer => d1_jtag_uart_0_avalon_jtag_slave_end_xfer,
      jtag_uart_0_avalon_jtag_slave_address => jtag_uart_0_avalon_jtag_slave_address,
      jtag_uart_0_avalon_jtag_slave_chipselect => jtag_uart_0_avalon_jtag_slave_chipselect,
      jtag_uart_0_avalon_jtag_slave_dataavailable_from_sa => jtag_uart_0_avalon_jtag_slave_dataavailable_from_sa,
      jtag_uart_0_avalon_jtag_slave_irq_from_sa => jtag_uart_0_avalon_jtag_slave_irq_from_sa,
      jtag_uart_0_avalon_jtag_slave_read_n => jtag_uart_0_avalon_jtag_slave_read_n,
      jtag_uart_0_avalon_jtag_slave_readdata_from_sa => jtag_uart_0_avalon_jtag_slave_readdata_from_sa,
      jtag_uart_0_avalon_jtag_slave_readyfordata_from_sa => jtag_uart_0_avalon_jtag_slave_readyfordata_from_sa,
      jtag_uart_0_avalon_jtag_slave_reset_n => jtag_uart_0_avalon_jtag_slave_reset_n,
      jtag_uart_0_avalon_jtag_slave_waitrequest_from_sa => jtag_uart_0_avalon_jtag_slave_waitrequest_from_sa,
      jtag_uart_0_avalon_jtag_slave_write_n => jtag_uart_0_avalon_jtag_slave_write_n,
      jtag_uart_0_avalon_jtag_slave_writedata => jtag_uart_0_avalon_jtag_slave_writedata,
      niosII_openMac_clock_0_out_granted_jtag_uart_0_avalon_jtag_slave => niosII_openMac_clock_0_out_granted_jtag_uart_0_avalon_jtag_slave,
      niosII_openMac_clock_0_out_qualified_request_jtag_uart_0_avalon_jtag_slave => niosII_openMac_clock_0_out_qualified_request_jtag_uart_0_avalon_jtag_slave,
      niosII_openMac_clock_0_out_read_data_valid_jtag_uart_0_avalon_jtag_slave => niosII_openMac_clock_0_out_read_data_valid_jtag_uart_0_avalon_jtag_slave,
      niosII_openMac_clock_0_out_requests_jtag_uart_0_avalon_jtag_slave => niosII_openMac_clock_0_out_requests_jtag_uart_0_avalon_jtag_slave,
      clk => internal_clk50Meg,
      jtag_uart_0_avalon_jtag_slave_dataavailable => jtag_uart_0_avalon_jtag_slave_dataavailable,
      jtag_uart_0_avalon_jtag_slave_irq => jtag_uart_0_avalon_jtag_slave_irq,
      jtag_uart_0_avalon_jtag_slave_readdata => jtag_uart_0_avalon_jtag_slave_readdata,
      jtag_uart_0_avalon_jtag_slave_readyfordata => jtag_uart_0_avalon_jtag_slave_readyfordata,
      jtag_uart_0_avalon_jtag_slave_waitrequest => jtag_uart_0_avalon_jtag_slave_waitrequest,
      niosII_openMac_clock_0_out_address_to_slave => niosII_openMac_clock_0_out_address_to_slave,
      niosII_openMac_clock_0_out_nativeaddress => niosII_openMac_clock_0_out_nativeaddress,
      niosII_openMac_clock_0_out_read => niosII_openMac_clock_0_out_read,
      niosII_openMac_clock_0_out_write => niosII_openMac_clock_0_out_write,
      niosII_openMac_clock_0_out_writedata => niosII_openMac_clock_0_out_writedata,
      reset_n => clk50Meg_reset_n
    );


  --the_jtag_uart_0, which is an e_ptf_instance
  the_jtag_uart_0 : jtag_uart_0
    port map(
      av_irq => jtag_uart_0_avalon_jtag_slave_irq,
      av_readdata => jtag_uart_0_avalon_jtag_slave_readdata,
      av_waitrequest => jtag_uart_0_avalon_jtag_slave_waitrequest,
      dataavailable => jtag_uart_0_avalon_jtag_slave_dataavailable,
      readyfordata => jtag_uart_0_avalon_jtag_slave_readyfordata,
      av_address => jtag_uart_0_avalon_jtag_slave_address,
      av_chipselect => jtag_uart_0_avalon_jtag_slave_chipselect,
      av_read_n => jtag_uart_0_avalon_jtag_slave_read_n,
      av_write_n => jtag_uart_0_avalon_jtag_slave_write_n,
      av_writedata => jtag_uart_0_avalon_jtag_slave_writedata,
      clk => internal_clk50Meg,
      rst_n => jtag_uart_0_avalon_jtag_slave_reset_n
    );


  --the_jtag_uart_1_avalon_jtag_slave, which is an e_instance
  the_jtag_uart_1_avalon_jtag_slave : jtag_uart_1_avalon_jtag_slave_arbitrator
    port map(
      ap_cpu_data_master_granted_jtag_uart_1_avalon_jtag_slave => ap_cpu_data_master_granted_jtag_uart_1_avalon_jtag_slave,
      ap_cpu_data_master_qualified_request_jtag_uart_1_avalon_jtag_slave => ap_cpu_data_master_qualified_request_jtag_uart_1_avalon_jtag_slave,
      ap_cpu_data_master_read_data_valid_jtag_uart_1_avalon_jtag_slave => ap_cpu_data_master_read_data_valid_jtag_uart_1_avalon_jtag_slave,
      ap_cpu_data_master_requests_jtag_uart_1_avalon_jtag_slave => ap_cpu_data_master_requests_jtag_uart_1_avalon_jtag_slave,
      d1_jtag_uart_1_avalon_jtag_slave_end_xfer => d1_jtag_uart_1_avalon_jtag_slave_end_xfer,
      jtag_uart_1_avalon_jtag_slave_address => jtag_uart_1_avalon_jtag_slave_address,
      jtag_uart_1_avalon_jtag_slave_chipselect => jtag_uart_1_avalon_jtag_slave_chipselect,
      jtag_uart_1_avalon_jtag_slave_dataavailable_from_sa => jtag_uart_1_avalon_jtag_slave_dataavailable_from_sa,
      jtag_uart_1_avalon_jtag_slave_irq_from_sa => jtag_uart_1_avalon_jtag_slave_irq_from_sa,
      jtag_uart_1_avalon_jtag_slave_read_n => jtag_uart_1_avalon_jtag_slave_read_n,
      jtag_uart_1_avalon_jtag_slave_readdata_from_sa => jtag_uart_1_avalon_jtag_slave_readdata_from_sa,
      jtag_uart_1_avalon_jtag_slave_readyfordata_from_sa => jtag_uart_1_avalon_jtag_slave_readyfordata_from_sa,
      jtag_uart_1_avalon_jtag_slave_reset_n => jtag_uart_1_avalon_jtag_slave_reset_n,
      jtag_uart_1_avalon_jtag_slave_waitrequest_from_sa => jtag_uart_1_avalon_jtag_slave_waitrequest_from_sa,
      jtag_uart_1_avalon_jtag_slave_write_n => jtag_uart_1_avalon_jtag_slave_write_n,
      jtag_uart_1_avalon_jtag_slave_writedata => jtag_uart_1_avalon_jtag_slave_writedata,
      ap_cpu_data_master_address_to_slave => ap_cpu_data_master_address_to_slave,
      ap_cpu_data_master_read => ap_cpu_data_master_read,
      ap_cpu_data_master_waitrequest => ap_cpu_data_master_waitrequest,
      ap_cpu_data_master_write => ap_cpu_data_master_write,
      ap_cpu_data_master_writedata => ap_cpu_data_master_writedata,
      clk => internal_clk90Meg,
      jtag_uart_1_avalon_jtag_slave_dataavailable => jtag_uart_1_avalon_jtag_slave_dataavailable,
      jtag_uart_1_avalon_jtag_slave_irq => jtag_uart_1_avalon_jtag_slave_irq,
      jtag_uart_1_avalon_jtag_slave_readdata => jtag_uart_1_avalon_jtag_slave_readdata,
      jtag_uart_1_avalon_jtag_slave_readyfordata => jtag_uart_1_avalon_jtag_slave_readyfordata,
      jtag_uart_1_avalon_jtag_slave_waitrequest => jtag_uart_1_avalon_jtag_slave_waitrequest,
      reset_n => clk90Meg_reset_n
    );


  --the_jtag_uart_1, which is an e_ptf_instance
  the_jtag_uart_1 : jtag_uart_1
    port map(
      av_irq => jtag_uart_1_avalon_jtag_slave_irq,
      av_readdata => jtag_uart_1_avalon_jtag_slave_readdata,
      av_waitrequest => jtag_uart_1_avalon_jtag_slave_waitrequest,
      dataavailable => jtag_uart_1_avalon_jtag_slave_dataavailable,
      readyfordata => jtag_uart_1_avalon_jtag_slave_readyfordata,
      av_address => jtag_uart_1_avalon_jtag_slave_address,
      av_chipselect => jtag_uart_1_avalon_jtag_slave_chipselect,
      av_read_n => jtag_uart_1_avalon_jtag_slave_read_n,
      av_write_n => jtag_uart_1_avalon_jtag_slave_write_n,
      av_writedata => jtag_uart_1_avalon_jtag_slave_writedata,
      clk => internal_clk90Meg,
      rst_n => jtag_uart_1_avalon_jtag_slave_reset_n
    );


  --the_niosII_openMac_clock_0_in, which is an e_instance
  the_niosII_openMac_clock_0_in : niosII_openMac_clock_0_in_arbitrator
    port map(
      d1_niosII_openMac_clock_0_in_end_xfer => d1_niosII_openMac_clock_0_in_end_xfer,
      niosII_openMac_clock_0_in_address => niosII_openMac_clock_0_in_address,
      niosII_openMac_clock_0_in_byteenable => niosII_openMac_clock_0_in_byteenable,
      niosII_openMac_clock_0_in_endofpacket_from_sa => niosII_openMac_clock_0_in_endofpacket_from_sa,
      niosII_openMac_clock_0_in_nativeaddress => niosII_openMac_clock_0_in_nativeaddress,
      niosII_openMac_clock_0_in_read => niosII_openMac_clock_0_in_read,
      niosII_openMac_clock_0_in_readdata_from_sa => niosII_openMac_clock_0_in_readdata_from_sa,
      niosII_openMac_clock_0_in_reset_n => niosII_openMac_clock_0_in_reset_n,
      niosII_openMac_clock_0_in_waitrequest_from_sa => niosII_openMac_clock_0_in_waitrequest_from_sa,
      niosII_openMac_clock_0_in_write => niosII_openMac_clock_0_in_write,
      niosII_openMac_clock_0_in_writedata => niosII_openMac_clock_0_in_writedata,
      pcp_cpu_data_master_granted_niosII_openMac_clock_0_in => pcp_cpu_data_master_granted_niosII_openMac_clock_0_in,
      pcp_cpu_data_master_qualified_request_niosII_openMac_clock_0_in => pcp_cpu_data_master_qualified_request_niosII_openMac_clock_0_in,
      pcp_cpu_data_master_read_data_valid_niosII_openMac_clock_0_in => pcp_cpu_data_master_read_data_valid_niosII_openMac_clock_0_in,
      pcp_cpu_data_master_requests_niosII_openMac_clock_0_in => pcp_cpu_data_master_requests_niosII_openMac_clock_0_in,
      clk => internal_clk90Meg,
      niosII_openMac_clock_0_in_endofpacket => niosII_openMac_clock_0_in_endofpacket,
      niosII_openMac_clock_0_in_readdata => niosII_openMac_clock_0_in_readdata,
      niosII_openMac_clock_0_in_waitrequest => niosII_openMac_clock_0_in_waitrequest,
      pcp_cpu_data_master_address_to_slave => pcp_cpu_data_master_address_to_slave,
      pcp_cpu_data_master_byteenable => pcp_cpu_data_master_byteenable,
      pcp_cpu_data_master_read => pcp_cpu_data_master_read,
      pcp_cpu_data_master_waitrequest => pcp_cpu_data_master_waitrequest,
      pcp_cpu_data_master_write => pcp_cpu_data_master_write,
      pcp_cpu_data_master_writedata => pcp_cpu_data_master_writedata,
      reset_n => clk90Meg_reset_n
    );


  --the_niosII_openMac_clock_0_out, which is an e_instance
  the_niosII_openMac_clock_0_out : niosII_openMac_clock_0_out_arbitrator
    port map(
      niosII_openMac_clock_0_out_address_to_slave => niosII_openMac_clock_0_out_address_to_slave,
      niosII_openMac_clock_0_out_readdata => niosII_openMac_clock_0_out_readdata,
      niosII_openMac_clock_0_out_reset_n => niosII_openMac_clock_0_out_reset_n,
      niosII_openMac_clock_0_out_waitrequest => niosII_openMac_clock_0_out_waitrequest,
      clk => internal_clk50Meg,
      d1_jtag_uart_0_avalon_jtag_slave_end_xfer => d1_jtag_uart_0_avalon_jtag_slave_end_xfer,
      jtag_uart_0_avalon_jtag_slave_readdata_from_sa => jtag_uart_0_avalon_jtag_slave_readdata_from_sa,
      jtag_uart_0_avalon_jtag_slave_waitrequest_from_sa => jtag_uart_0_avalon_jtag_slave_waitrequest_from_sa,
      niosII_openMac_clock_0_out_address => niosII_openMac_clock_0_out_address,
      niosII_openMac_clock_0_out_byteenable => niosII_openMac_clock_0_out_byteenable,
      niosII_openMac_clock_0_out_granted_jtag_uart_0_avalon_jtag_slave => niosII_openMac_clock_0_out_granted_jtag_uart_0_avalon_jtag_slave,
      niosII_openMac_clock_0_out_qualified_request_jtag_uart_0_avalon_jtag_slave => niosII_openMac_clock_0_out_qualified_request_jtag_uart_0_avalon_jtag_slave,
      niosII_openMac_clock_0_out_read => niosII_openMac_clock_0_out_read,
      niosII_openMac_clock_0_out_read_data_valid_jtag_uart_0_avalon_jtag_slave => niosII_openMac_clock_0_out_read_data_valid_jtag_uart_0_avalon_jtag_slave,
      niosII_openMac_clock_0_out_requests_jtag_uart_0_avalon_jtag_slave => niosII_openMac_clock_0_out_requests_jtag_uart_0_avalon_jtag_slave,
      niosII_openMac_clock_0_out_write => niosII_openMac_clock_0_out_write,
      niosII_openMac_clock_0_out_writedata => niosII_openMac_clock_0_out_writedata,
      reset_n => clk50Meg_reset_n
    );


  --the_niosII_openMac_clock_0, which is an e_ptf_instance
  the_niosII_openMac_clock_0 : niosII_openMac_clock_0
    port map(
      master_address => niosII_openMac_clock_0_out_address,
      master_byteenable => niosII_openMac_clock_0_out_byteenable,
      master_nativeaddress => niosII_openMac_clock_0_out_nativeaddress,
      master_read => niosII_openMac_clock_0_out_read,
      master_write => niosII_openMac_clock_0_out_write,
      master_writedata => niosII_openMac_clock_0_out_writedata,
      slave_endofpacket => niosII_openMac_clock_0_in_endofpacket,
      slave_readdata => niosII_openMac_clock_0_in_readdata,
      slave_waitrequest => niosII_openMac_clock_0_in_waitrequest,
      master_clk => internal_clk50Meg,
      master_endofpacket => niosII_openMac_clock_0_out_endofpacket,
      master_readdata => niosII_openMac_clock_0_out_readdata,
      master_reset_n => niosII_openMac_clock_0_out_reset_n,
      master_waitrequest => niosII_openMac_clock_0_out_waitrequest,
      slave_address => niosII_openMac_clock_0_in_address,
      slave_byteenable => niosII_openMac_clock_0_in_byteenable,
      slave_clk => internal_clk90Meg,
      slave_nativeaddress => niosII_openMac_clock_0_in_nativeaddress,
      slave_read => niosII_openMac_clock_0_in_read,
      slave_reset_n => niosII_openMac_clock_0_in_reset_n,
      slave_write => niosII_openMac_clock_0_in_write,
      slave_writedata => niosII_openMac_clock_0_in_writedata
    );


  --the_niosII_openMac_clock_1_in, which is an e_instance
  the_niosII_openMac_clock_1_in : niosII_openMac_clock_1_in_arbitrator
    port map(
      d1_niosII_openMac_clock_1_in_end_xfer => d1_niosII_openMac_clock_1_in_end_xfer,
      niosII_openMac_clock_1_in_address => niosII_openMac_clock_1_in_address,
      niosII_openMac_clock_1_in_byteenable => niosII_openMac_clock_1_in_byteenable,
      niosII_openMac_clock_1_in_endofpacket_from_sa => niosII_openMac_clock_1_in_endofpacket_from_sa,
      niosII_openMac_clock_1_in_nativeaddress => niosII_openMac_clock_1_in_nativeaddress,
      niosII_openMac_clock_1_in_read => niosII_openMac_clock_1_in_read,
      niosII_openMac_clock_1_in_readdata_from_sa => niosII_openMac_clock_1_in_readdata_from_sa,
      niosII_openMac_clock_1_in_reset_n => niosII_openMac_clock_1_in_reset_n,
      niosII_openMac_clock_1_in_waitrequest_from_sa => niosII_openMac_clock_1_in_waitrequest_from_sa,
      niosII_openMac_clock_1_in_write => niosII_openMac_clock_1_in_write,
      niosII_openMac_clock_1_in_writedata => niosII_openMac_clock_1_in_writedata,
      pcp_cpu_data_master_granted_niosII_openMac_clock_1_in => pcp_cpu_data_master_granted_niosII_openMac_clock_1_in,
      pcp_cpu_data_master_qualified_request_niosII_openMac_clock_1_in => pcp_cpu_data_master_qualified_request_niosII_openMac_clock_1_in,
      pcp_cpu_data_master_read_data_valid_niosII_openMac_clock_1_in => pcp_cpu_data_master_read_data_valid_niosII_openMac_clock_1_in,
      pcp_cpu_data_master_requests_niosII_openMac_clock_1_in => pcp_cpu_data_master_requests_niosII_openMac_clock_1_in,
      clk => internal_clk90Meg,
      niosII_openMac_clock_1_in_endofpacket => niosII_openMac_clock_1_in_endofpacket,
      niosII_openMac_clock_1_in_readdata => niosII_openMac_clock_1_in_readdata,
      niosII_openMac_clock_1_in_waitrequest => niosII_openMac_clock_1_in_waitrequest,
      pcp_cpu_data_master_address_to_slave => pcp_cpu_data_master_address_to_slave,
      pcp_cpu_data_master_byteenable => pcp_cpu_data_master_byteenable,
      pcp_cpu_data_master_read => pcp_cpu_data_master_read,
      pcp_cpu_data_master_waitrequest => pcp_cpu_data_master_waitrequest,
      pcp_cpu_data_master_write => pcp_cpu_data_master_write,
      pcp_cpu_data_master_writedata => pcp_cpu_data_master_writedata,
      reset_n => clk90Meg_reset_n
    );


  --the_niosII_openMac_clock_1_out, which is an e_instance
  the_niosII_openMac_clock_1_out : niosII_openMac_clock_1_out_arbitrator
    port map(
      niosII_openMac_clock_1_out_address_to_slave => niosII_openMac_clock_1_out_address_to_slave,
      niosII_openMac_clock_1_out_readdata => niosII_openMac_clock_1_out_readdata,
      niosII_openMac_clock_1_out_reset_n => niosII_openMac_clock_1_out_reset_n,
      niosII_openMac_clock_1_out_waitrequest => niosII_openMac_clock_1_out_waitrequest,
      OpenMAC_0_CMP_readdata_from_sa => OpenMAC_0_CMP_readdata_from_sa,
      clk => internal_clk50Meg,
      d1_OpenMAC_0_CMP_end_xfer => d1_OpenMAC_0_CMP_end_xfer,
      niosII_openMac_clock_1_out_address => niosII_openMac_clock_1_out_address,
      niosII_openMac_clock_1_out_byteenable => niosII_openMac_clock_1_out_byteenable,
      niosII_openMac_clock_1_out_granted_OpenMAC_0_CMP => niosII_openMac_clock_1_out_granted_OpenMAC_0_CMP,
      niosII_openMac_clock_1_out_qualified_request_OpenMAC_0_CMP => niosII_openMac_clock_1_out_qualified_request_OpenMAC_0_CMP,
      niosII_openMac_clock_1_out_read => niosII_openMac_clock_1_out_read,
      niosII_openMac_clock_1_out_read_data_valid_OpenMAC_0_CMP => niosII_openMac_clock_1_out_read_data_valid_OpenMAC_0_CMP,
      niosII_openMac_clock_1_out_requests_OpenMAC_0_CMP => niosII_openMac_clock_1_out_requests_OpenMAC_0_CMP,
      niosII_openMac_clock_1_out_write => niosII_openMac_clock_1_out_write,
      niosII_openMac_clock_1_out_writedata => niosII_openMac_clock_1_out_writedata,
      reset_n => clk50Meg_reset_n
    );


  --the_niosII_openMac_clock_1, which is an e_ptf_instance
  the_niosII_openMac_clock_1 : niosII_openMac_clock_1
    port map(
      master_address => niosII_openMac_clock_1_out_address,
      master_byteenable => niosII_openMac_clock_1_out_byteenable,
      master_nativeaddress => niosII_openMac_clock_1_out_nativeaddress,
      master_read => niosII_openMac_clock_1_out_read,
      master_write => niosII_openMac_clock_1_out_write,
      master_writedata => niosII_openMac_clock_1_out_writedata,
      slave_endofpacket => niosII_openMac_clock_1_in_endofpacket,
      slave_readdata => niosII_openMac_clock_1_in_readdata,
      slave_waitrequest => niosII_openMac_clock_1_in_waitrequest,
      master_clk => internal_clk50Meg,
      master_endofpacket => niosII_openMac_clock_1_out_endofpacket,
      master_readdata => niosII_openMac_clock_1_out_readdata,
      master_reset_n => niosII_openMac_clock_1_out_reset_n,
      master_waitrequest => niosII_openMac_clock_1_out_waitrequest,
      slave_address => niosII_openMac_clock_1_in_address,
      slave_byteenable => niosII_openMac_clock_1_in_byteenable,
      slave_clk => internal_clk90Meg,
      slave_nativeaddress => niosII_openMac_clock_1_in_nativeaddress,
      slave_read => niosII_openMac_clock_1_in_read,
      slave_reset_n => niosII_openMac_clock_1_in_reset_n,
      slave_write => niosII_openMac_clock_1_in_write,
      slave_writedata => niosII_openMac_clock_1_in_writedata
    );


  --the_niosII_openMac_clock_2_in, which is an e_instance
  the_niosII_openMac_clock_2_in : niosII_openMac_clock_2_in_arbitrator
    port map(
      d1_niosII_openMac_clock_2_in_end_xfer => d1_niosII_openMac_clock_2_in_end_xfer,
      niosII_openMac_clock_2_in_address => niosII_openMac_clock_2_in_address,
      niosII_openMac_clock_2_in_byteenable => niosII_openMac_clock_2_in_byteenable,
      niosII_openMac_clock_2_in_endofpacket_from_sa => niosII_openMac_clock_2_in_endofpacket_from_sa,
      niosII_openMac_clock_2_in_nativeaddress => niosII_openMac_clock_2_in_nativeaddress,
      niosII_openMac_clock_2_in_read => niosII_openMac_clock_2_in_read,
      niosII_openMac_clock_2_in_readdata_from_sa => niosII_openMac_clock_2_in_readdata_from_sa,
      niosII_openMac_clock_2_in_reset_n => niosII_openMac_clock_2_in_reset_n,
      niosII_openMac_clock_2_in_waitrequest_from_sa => niosII_openMac_clock_2_in_waitrequest_from_sa,
      niosII_openMac_clock_2_in_write => niosII_openMac_clock_2_in_write,
      niosII_openMac_clock_2_in_writedata => niosII_openMac_clock_2_in_writedata,
      pcp_cpu_data_master_byteenable_niosII_openMac_clock_2_in => pcp_cpu_data_master_byteenable_niosII_openMac_clock_2_in,
      pcp_cpu_data_master_granted_niosII_openMac_clock_2_in => pcp_cpu_data_master_granted_niosII_openMac_clock_2_in,
      pcp_cpu_data_master_qualified_request_niosII_openMac_clock_2_in => pcp_cpu_data_master_qualified_request_niosII_openMac_clock_2_in,
      pcp_cpu_data_master_read_data_valid_niosII_openMac_clock_2_in => pcp_cpu_data_master_read_data_valid_niosII_openMac_clock_2_in,
      pcp_cpu_data_master_requests_niosII_openMac_clock_2_in => pcp_cpu_data_master_requests_niosII_openMac_clock_2_in,
      clk => internal_clk90Meg,
      niosII_openMac_clock_2_in_endofpacket => niosII_openMac_clock_2_in_endofpacket,
      niosII_openMac_clock_2_in_readdata => niosII_openMac_clock_2_in_readdata,
      niosII_openMac_clock_2_in_waitrequest => niosII_openMac_clock_2_in_waitrequest,
      pcp_cpu_data_master_address_to_slave => pcp_cpu_data_master_address_to_slave,
      pcp_cpu_data_master_byteenable => pcp_cpu_data_master_byteenable,
      pcp_cpu_data_master_dbs_address => pcp_cpu_data_master_dbs_address,
      pcp_cpu_data_master_dbs_write_16 => pcp_cpu_data_master_dbs_write_16,
      pcp_cpu_data_master_no_byte_enables_and_last_term => pcp_cpu_data_master_no_byte_enables_and_last_term,
      pcp_cpu_data_master_read => pcp_cpu_data_master_read,
      pcp_cpu_data_master_waitrequest => pcp_cpu_data_master_waitrequest,
      pcp_cpu_data_master_write => pcp_cpu_data_master_write,
      reset_n => clk90Meg_reset_n
    );


  --the_niosII_openMac_clock_2_out, which is an e_instance
  the_niosII_openMac_clock_2_out : niosII_openMac_clock_2_out_arbitrator
    port map(
      niosII_openMac_clock_2_out_address_to_slave => niosII_openMac_clock_2_out_address_to_slave,
      niosII_openMac_clock_2_out_readdata => niosII_openMac_clock_2_out_readdata,
      niosII_openMac_clock_2_out_reset_n => niosII_openMac_clock_2_out_reset_n,
      niosII_openMac_clock_2_out_waitrequest => niosII_openMac_clock_2_out_waitrequest,
      OpenMAC_0_REG_readdata_from_sa => OpenMAC_0_REG_readdata_from_sa,
      clk => internal_clk50Meg,
      d1_OpenMAC_0_REG_end_xfer => d1_OpenMAC_0_REG_end_xfer,
      niosII_openMac_clock_2_out_address => niosII_openMac_clock_2_out_address,
      niosII_openMac_clock_2_out_byteenable => niosII_openMac_clock_2_out_byteenable,
      niosII_openMac_clock_2_out_granted_OpenMAC_0_REG => niosII_openMac_clock_2_out_granted_OpenMAC_0_REG,
      niosII_openMac_clock_2_out_qualified_request_OpenMAC_0_REG => niosII_openMac_clock_2_out_qualified_request_OpenMAC_0_REG,
      niosII_openMac_clock_2_out_read => niosII_openMac_clock_2_out_read,
      niosII_openMac_clock_2_out_read_data_valid_OpenMAC_0_REG => niosII_openMac_clock_2_out_read_data_valid_OpenMAC_0_REG,
      niosII_openMac_clock_2_out_requests_OpenMAC_0_REG => niosII_openMac_clock_2_out_requests_OpenMAC_0_REG,
      niosII_openMac_clock_2_out_write => niosII_openMac_clock_2_out_write,
      niosII_openMac_clock_2_out_writedata => niosII_openMac_clock_2_out_writedata,
      reset_n => clk50Meg_reset_n
    );


  --the_niosII_openMac_clock_2, which is an e_ptf_instance
  the_niosII_openMac_clock_2 : niosII_openMac_clock_2
    port map(
      master_address => niosII_openMac_clock_2_out_address,
      master_byteenable => niosII_openMac_clock_2_out_byteenable,
      master_nativeaddress => niosII_openMac_clock_2_out_nativeaddress,
      master_read => niosII_openMac_clock_2_out_read,
      master_write => niosII_openMac_clock_2_out_write,
      master_writedata => niosII_openMac_clock_2_out_writedata,
      slave_endofpacket => niosII_openMac_clock_2_in_endofpacket,
      slave_readdata => niosII_openMac_clock_2_in_readdata,
      slave_waitrequest => niosII_openMac_clock_2_in_waitrequest,
      master_clk => internal_clk50Meg,
      master_endofpacket => niosII_openMac_clock_2_out_endofpacket,
      master_readdata => niosII_openMac_clock_2_out_readdata,
      master_reset_n => niosII_openMac_clock_2_out_reset_n,
      master_waitrequest => niosII_openMac_clock_2_out_waitrequest,
      slave_address => niosII_openMac_clock_2_in_address,
      slave_byteenable => niosII_openMac_clock_2_in_byteenable,
      slave_clk => internal_clk90Meg,
      slave_nativeaddress => niosII_openMac_clock_2_in_nativeaddress,
      slave_read => niosII_openMac_clock_2_in_read,
      slave_reset_n => niosII_openMac_clock_2_in_reset_n,
      slave_write => niosII_openMac_clock_2_in_write,
      slave_writedata => niosII_openMac_clock_2_in_writedata
    );


  --the_niosII_openMac_clock_3_in, which is an e_instance
  the_niosII_openMac_clock_3_in : niosII_openMac_clock_3_in_arbitrator
    port map(
      d1_niosII_openMac_clock_3_in_end_xfer => d1_niosII_openMac_clock_3_in_end_xfer,
      niosII_openMac_clock_3_in_address => niosII_openMac_clock_3_in_address,
      niosII_openMac_clock_3_in_byteenable => niosII_openMac_clock_3_in_byteenable,
      niosII_openMac_clock_3_in_endofpacket_from_sa => niosII_openMac_clock_3_in_endofpacket_from_sa,
      niosII_openMac_clock_3_in_nativeaddress => niosII_openMac_clock_3_in_nativeaddress,
      niosII_openMac_clock_3_in_read => niosII_openMac_clock_3_in_read,
      niosII_openMac_clock_3_in_readdata_from_sa => niosII_openMac_clock_3_in_readdata_from_sa,
      niosII_openMac_clock_3_in_reset_n => niosII_openMac_clock_3_in_reset_n,
      niosII_openMac_clock_3_in_waitrequest_from_sa => niosII_openMac_clock_3_in_waitrequest_from_sa,
      niosII_openMac_clock_3_in_write => niosII_openMac_clock_3_in_write,
      niosII_openMac_clock_3_in_writedata => niosII_openMac_clock_3_in_writedata,
      pcp_cpu_data_master_granted_niosII_openMac_clock_3_in => pcp_cpu_data_master_granted_niosII_openMac_clock_3_in,
      pcp_cpu_data_master_qualified_request_niosII_openMac_clock_3_in => pcp_cpu_data_master_qualified_request_niosII_openMac_clock_3_in,
      pcp_cpu_data_master_read_data_valid_niosII_openMac_clock_3_in => pcp_cpu_data_master_read_data_valid_niosII_openMac_clock_3_in,
      pcp_cpu_data_master_requests_niosII_openMac_clock_3_in => pcp_cpu_data_master_requests_niosII_openMac_clock_3_in,
      clk => internal_clk90Meg,
      niosII_openMac_clock_3_in_endofpacket => niosII_openMac_clock_3_in_endofpacket,
      niosII_openMac_clock_3_in_readdata => niosII_openMac_clock_3_in_readdata,
      niosII_openMac_clock_3_in_waitrequest => niosII_openMac_clock_3_in_waitrequest,
      pcp_cpu_data_master_address_to_slave => pcp_cpu_data_master_address_to_slave,
      pcp_cpu_data_master_byteenable => pcp_cpu_data_master_byteenable,
      pcp_cpu_data_master_read => pcp_cpu_data_master_read,
      pcp_cpu_data_master_waitrequest => pcp_cpu_data_master_waitrequest,
      pcp_cpu_data_master_write => pcp_cpu_data_master_write,
      pcp_cpu_data_master_writedata => pcp_cpu_data_master_writedata,
      reset_n => clk90Meg_reset_n
    );


  --the_niosII_openMac_clock_3_out, which is an e_instance
  the_niosII_openMac_clock_3_out : niosII_openMac_clock_3_out_arbitrator
    port map(
      niosII_openMac_clock_3_out_address_to_slave => niosII_openMac_clock_3_out_address_to_slave,
      niosII_openMac_clock_3_out_readdata => niosII_openMac_clock_3_out_readdata,
      niosII_openMac_clock_3_out_reset_n => niosII_openMac_clock_3_out_reset_n,
      niosII_openMac_clock_3_out_waitrequest => niosII_openMac_clock_3_out_waitrequest,
      altpll_0_pll_slave_readdata_from_sa => altpll_0_pll_slave_readdata_from_sa,
      clk => clk_0,
      d1_altpll_0_pll_slave_end_xfer => d1_altpll_0_pll_slave_end_xfer,
      niosII_openMac_clock_3_out_address => niosII_openMac_clock_3_out_address,
      niosII_openMac_clock_3_out_byteenable => niosII_openMac_clock_3_out_byteenable,
      niosII_openMac_clock_3_out_granted_altpll_0_pll_slave => niosII_openMac_clock_3_out_granted_altpll_0_pll_slave,
      niosII_openMac_clock_3_out_qualified_request_altpll_0_pll_slave => niosII_openMac_clock_3_out_qualified_request_altpll_0_pll_slave,
      niosII_openMac_clock_3_out_read => niosII_openMac_clock_3_out_read,
      niosII_openMac_clock_3_out_read_data_valid_altpll_0_pll_slave => niosII_openMac_clock_3_out_read_data_valid_altpll_0_pll_slave,
      niosII_openMac_clock_3_out_requests_altpll_0_pll_slave => niosII_openMac_clock_3_out_requests_altpll_0_pll_slave,
      niosII_openMac_clock_3_out_write => niosII_openMac_clock_3_out_write,
      niosII_openMac_clock_3_out_writedata => niosII_openMac_clock_3_out_writedata,
      reset_n => clk_0_reset_n
    );


  --the_niosII_openMac_clock_3, which is an e_ptf_instance
  the_niosII_openMac_clock_3 : niosII_openMac_clock_3
    port map(
      master_address => niosII_openMac_clock_3_out_address,
      master_byteenable => niosII_openMac_clock_3_out_byteenable,
      master_nativeaddress => niosII_openMac_clock_3_out_nativeaddress,
      master_read => niosII_openMac_clock_3_out_read,
      master_write => niosII_openMac_clock_3_out_write,
      master_writedata => niosII_openMac_clock_3_out_writedata,
      slave_endofpacket => niosII_openMac_clock_3_in_endofpacket,
      slave_readdata => niosII_openMac_clock_3_in_readdata,
      slave_waitrequest => niosII_openMac_clock_3_in_waitrequest,
      master_clk => clk_0,
      master_endofpacket => niosII_openMac_clock_3_out_endofpacket,
      master_readdata => niosII_openMac_clock_3_out_readdata,
      master_reset_n => niosII_openMac_clock_3_out_reset_n,
      master_waitrequest => niosII_openMac_clock_3_out_waitrequest,
      slave_address => niosII_openMac_clock_3_in_address,
      slave_byteenable => niosII_openMac_clock_3_in_byteenable,
      slave_clk => internal_clk90Meg,
      slave_nativeaddress => niosII_openMac_clock_3_in_nativeaddress,
      slave_read => niosII_openMac_clock_3_in_read,
      slave_reset_n => niosII_openMac_clock_3_in_reset_n,
      slave_write => niosII_openMac_clock_3_in_write,
      slave_writedata => niosII_openMac_clock_3_in_writedata
    );


  --the_niosII_openMac_clock_4_in, which is an e_instance
  the_niosII_openMac_clock_4_in : niosII_openMac_clock_4_in_arbitrator
    port map(
      d1_niosII_openMac_clock_4_in_end_xfer => d1_niosII_openMac_clock_4_in_end_xfer,
      niosII_openMac_clock_4_in_address => niosII_openMac_clock_4_in_address,
      niosII_openMac_clock_4_in_byteenable => niosII_openMac_clock_4_in_byteenable,
      niosII_openMac_clock_4_in_endofpacket_from_sa => niosII_openMac_clock_4_in_endofpacket_from_sa,
      niosII_openMac_clock_4_in_nativeaddress => niosII_openMac_clock_4_in_nativeaddress,
      niosII_openMac_clock_4_in_read => niosII_openMac_clock_4_in_read,
      niosII_openMac_clock_4_in_readdata_from_sa => niosII_openMac_clock_4_in_readdata_from_sa,
      niosII_openMac_clock_4_in_reset_n => niosII_openMac_clock_4_in_reset_n,
      niosII_openMac_clock_4_in_waitrequest_from_sa => niosII_openMac_clock_4_in_waitrequest_from_sa,
      niosII_openMac_clock_4_in_write => niosII_openMac_clock_4_in_write,
      niosII_openMac_clock_4_in_writedata => niosII_openMac_clock_4_in_writedata,
      pcp_cpu_data_master_granted_niosII_openMac_clock_4_in => pcp_cpu_data_master_granted_niosII_openMac_clock_4_in,
      pcp_cpu_data_master_qualified_request_niosII_openMac_clock_4_in => pcp_cpu_data_master_qualified_request_niosII_openMac_clock_4_in,
      pcp_cpu_data_master_read_data_valid_niosII_openMac_clock_4_in => pcp_cpu_data_master_read_data_valid_niosII_openMac_clock_4_in,
      pcp_cpu_data_master_requests_niosII_openMac_clock_4_in => pcp_cpu_data_master_requests_niosII_openMac_clock_4_in,
      clk => internal_clk90Meg,
      niosII_openMac_clock_4_in_endofpacket => niosII_openMac_clock_4_in_endofpacket,
      niosII_openMac_clock_4_in_readdata => niosII_openMac_clock_4_in_readdata,
      niosII_openMac_clock_4_in_waitrequest => niosII_openMac_clock_4_in_waitrequest,
      pcp_cpu_data_master_address_to_slave => pcp_cpu_data_master_address_to_slave,
      pcp_cpu_data_master_byteenable => pcp_cpu_data_master_byteenable,
      pcp_cpu_data_master_read => pcp_cpu_data_master_read,
      pcp_cpu_data_master_waitrequest => pcp_cpu_data_master_waitrequest,
      pcp_cpu_data_master_write => pcp_cpu_data_master_write,
      pcp_cpu_data_master_writedata => pcp_cpu_data_master_writedata,
      reset_n => clk90Meg_reset_n
    );


  --the_niosII_openMac_clock_4_out, which is an e_instance
  the_niosII_openMac_clock_4_out : niosII_openMac_clock_4_out_arbitrator
    port map(
      niosII_openMac_clock_4_out_address_to_slave => niosII_openMac_clock_4_out_address_to_slave,
      niosII_openMac_clock_4_out_readdata => niosII_openMac_clock_4_out_readdata,
      niosII_openMac_clock_4_out_reset_n => niosII_openMac_clock_4_out_reset_n,
      niosII_openMac_clock_4_out_waitrequest => niosII_openMac_clock_4_out_waitrequest,
      clk => internal_clk25Meg,
      d1_remote_update_cycloneiii_0_s1_end_xfer => d1_remote_update_cycloneiii_0_s1_end_xfer,
      niosII_openMac_clock_4_out_address => niosII_openMac_clock_4_out_address,
      niosII_openMac_clock_4_out_byteenable => niosII_openMac_clock_4_out_byteenable,
      niosII_openMac_clock_4_out_granted_remote_update_cycloneiii_0_s1 => niosII_openMac_clock_4_out_granted_remote_update_cycloneiii_0_s1,
      niosII_openMac_clock_4_out_qualified_request_remote_update_cycloneiii_0_s1 => niosII_openMac_clock_4_out_qualified_request_remote_update_cycloneiii_0_s1,
      niosII_openMac_clock_4_out_read => niosII_openMac_clock_4_out_read,
      niosII_openMac_clock_4_out_read_data_valid_remote_update_cycloneiii_0_s1 => niosII_openMac_clock_4_out_read_data_valid_remote_update_cycloneiii_0_s1,
      niosII_openMac_clock_4_out_requests_remote_update_cycloneiii_0_s1 => niosII_openMac_clock_4_out_requests_remote_update_cycloneiii_0_s1,
      niosII_openMac_clock_4_out_write => niosII_openMac_clock_4_out_write,
      niosII_openMac_clock_4_out_writedata => niosII_openMac_clock_4_out_writedata,
      remote_update_cycloneiii_0_s1_readdata_from_sa => remote_update_cycloneiii_0_s1_readdata_from_sa,
      remote_update_cycloneiii_0_s1_waitrequest_from_sa => remote_update_cycloneiii_0_s1_waitrequest_from_sa,
      reset_n => clk25Meg_reset_n
    );


  --the_niosII_openMac_clock_4, which is an e_ptf_instance
  the_niosII_openMac_clock_4 : niosII_openMac_clock_4
    port map(
      master_address => niosII_openMac_clock_4_out_address,
      master_byteenable => niosII_openMac_clock_4_out_byteenable,
      master_nativeaddress => niosII_openMac_clock_4_out_nativeaddress,
      master_read => niosII_openMac_clock_4_out_read,
      master_write => niosII_openMac_clock_4_out_write,
      master_writedata => niosII_openMac_clock_4_out_writedata,
      slave_endofpacket => niosII_openMac_clock_4_in_endofpacket,
      slave_readdata => niosII_openMac_clock_4_in_readdata,
      slave_waitrequest => niosII_openMac_clock_4_in_waitrequest,
      master_clk => internal_clk25Meg,
      master_endofpacket => niosII_openMac_clock_4_out_endofpacket,
      master_readdata => niosII_openMac_clock_4_out_readdata,
      master_reset_n => niosII_openMac_clock_4_out_reset_n,
      master_waitrequest => niosII_openMac_clock_4_out_waitrequest,
      slave_address => niosII_openMac_clock_4_in_address,
      slave_byteenable => niosII_openMac_clock_4_in_byteenable,
      slave_clk => internal_clk90Meg,
      slave_nativeaddress => niosII_openMac_clock_4_in_nativeaddress,
      slave_read => niosII_openMac_clock_4_in_read,
      slave_reset_n => niosII_openMac_clock_4_in_reset_n,
      slave_write => niosII_openMac_clock_4_in_write,
      slave_writedata => niosII_openMac_clock_4_in_writedata
    );


  --the_node_switch_pio_s1, which is an e_instance
  the_node_switch_pio_s1 : node_switch_pio_s1_arbitrator
    port map(
      clock_crossing_1_m1_granted_node_switch_pio_s1 => clock_crossing_1_m1_granted_node_switch_pio_s1,
      clock_crossing_1_m1_qualified_request_node_switch_pio_s1 => clock_crossing_1_m1_qualified_request_node_switch_pio_s1,
      clock_crossing_1_m1_read_data_valid_node_switch_pio_s1 => clock_crossing_1_m1_read_data_valid_node_switch_pio_s1,
      clock_crossing_1_m1_requests_node_switch_pio_s1 => clock_crossing_1_m1_requests_node_switch_pio_s1,
      d1_node_switch_pio_s1_end_xfer => d1_node_switch_pio_s1_end_xfer,
      node_switch_pio_s1_address => node_switch_pio_s1_address,
      node_switch_pio_s1_readdata_from_sa => node_switch_pio_s1_readdata_from_sa,
      node_switch_pio_s1_reset_n => node_switch_pio_s1_reset_n,
      clk => internal_clk50Meg,
      clock_crossing_1_m1_address_to_slave => clock_crossing_1_m1_address_to_slave,
      clock_crossing_1_m1_latency_counter => clock_crossing_1_m1_latency_counter,
      clock_crossing_1_m1_nativeaddress => clock_crossing_1_m1_nativeaddress,
      clock_crossing_1_m1_read => clock_crossing_1_m1_read,
      clock_crossing_1_m1_write => clock_crossing_1_m1_write,
      node_switch_pio_s1_readdata => node_switch_pio_s1_readdata,
      reset_n => clk50Meg_reset_n
    );


  --the_node_switch_pio, which is an e_ptf_instance
  the_node_switch_pio : node_switch_pio
    port map(
      readdata => node_switch_pio_s1_readdata,
      address => node_switch_pio_s1_address,
      clk => internal_clk50Meg,
      in_port => in_port_to_the_node_switch_pio,
      reset_n => node_switch_pio_s1_reset_n
    );


  --the_onchip_memory_0_s1, which is an e_instance
  the_onchip_memory_0_s1 : onchip_memory_0_s1_arbitrator
    port map(
      d1_onchip_memory_0_s1_end_xfer => d1_onchip_memory_0_s1_end_xfer,
      onchip_memory_0_s1_address => onchip_memory_0_s1_address,
      onchip_memory_0_s1_byteenable => onchip_memory_0_s1_byteenable,
      onchip_memory_0_s1_chipselect => onchip_memory_0_s1_chipselect,
      onchip_memory_0_s1_clken => onchip_memory_0_s1_clken,
      onchip_memory_0_s1_readdata_from_sa => onchip_memory_0_s1_readdata_from_sa,
      onchip_memory_0_s1_write => onchip_memory_0_s1_write,
      onchip_memory_0_s1_writedata => onchip_memory_0_s1_writedata,
      pcp_cpu_data_master_granted_onchip_memory_0_s1 => pcp_cpu_data_master_granted_onchip_memory_0_s1,
      pcp_cpu_data_master_qualified_request_onchip_memory_0_s1 => pcp_cpu_data_master_qualified_request_onchip_memory_0_s1,
      pcp_cpu_data_master_read_data_valid_onchip_memory_0_s1 => pcp_cpu_data_master_read_data_valid_onchip_memory_0_s1,
      pcp_cpu_data_master_requests_onchip_memory_0_s1 => pcp_cpu_data_master_requests_onchip_memory_0_s1,
      pcp_cpu_instruction_master_granted_onchip_memory_0_s1 => pcp_cpu_instruction_master_granted_onchip_memory_0_s1,
      pcp_cpu_instruction_master_qualified_request_onchip_memory_0_s1 => pcp_cpu_instruction_master_qualified_request_onchip_memory_0_s1,
      pcp_cpu_instruction_master_read_data_valid_onchip_memory_0_s1 => pcp_cpu_instruction_master_read_data_valid_onchip_memory_0_s1,
      pcp_cpu_instruction_master_requests_onchip_memory_0_s1 => pcp_cpu_instruction_master_requests_onchip_memory_0_s1,
      registered_pcp_cpu_data_master_read_data_valid_onchip_memory_0_s1 => registered_pcp_cpu_data_master_read_data_valid_onchip_memory_0_s1,
      clk => internal_clk90Meg,
      onchip_memory_0_s1_readdata => onchip_memory_0_s1_readdata,
      pcp_cpu_data_master_address_to_slave => pcp_cpu_data_master_address_to_slave,
      pcp_cpu_data_master_byteenable => pcp_cpu_data_master_byteenable,
      pcp_cpu_data_master_read => pcp_cpu_data_master_read,
      pcp_cpu_data_master_waitrequest => pcp_cpu_data_master_waitrequest,
      pcp_cpu_data_master_write => pcp_cpu_data_master_write,
      pcp_cpu_data_master_writedata => pcp_cpu_data_master_writedata,
      pcp_cpu_instruction_master_address_to_slave => pcp_cpu_instruction_master_address_to_slave,
      pcp_cpu_instruction_master_latency_counter => pcp_cpu_instruction_master_latency_counter,
      pcp_cpu_instruction_master_read => pcp_cpu_instruction_master_read,
      reset_n => clk90Meg_reset_n
    );


  --the_onchip_memory_0, which is an e_ptf_instance
  the_onchip_memory_0 : onchip_memory_0
    port map(
      readdata => onchip_memory_0_s1_readdata,
      address => onchip_memory_0_s1_address,
      byteenable => onchip_memory_0_s1_byteenable,
      chipselect => onchip_memory_0_s1_chipselect,
      clk => internal_clk90Meg,
      clken => onchip_memory_0_s1_clken,
      write => onchip_memory_0_s1_write,
      writedata => onchip_memory_0_s1_writedata
    );


  --the_pcp_cpu_jtag_debug_module, which is an e_instance
  the_pcp_cpu_jtag_debug_module : pcp_cpu_jtag_debug_module_arbitrator
    port map(
      d1_pcp_cpu_jtag_debug_module_end_xfer => d1_pcp_cpu_jtag_debug_module_end_xfer,
      pcp_cpu_data_master_granted_pcp_cpu_jtag_debug_module => pcp_cpu_data_master_granted_pcp_cpu_jtag_debug_module,
      pcp_cpu_data_master_qualified_request_pcp_cpu_jtag_debug_module => pcp_cpu_data_master_qualified_request_pcp_cpu_jtag_debug_module,
      pcp_cpu_data_master_read_data_valid_pcp_cpu_jtag_debug_module => pcp_cpu_data_master_read_data_valid_pcp_cpu_jtag_debug_module,
      pcp_cpu_data_master_requests_pcp_cpu_jtag_debug_module => pcp_cpu_data_master_requests_pcp_cpu_jtag_debug_module,
      pcp_cpu_instruction_master_granted_pcp_cpu_jtag_debug_module => pcp_cpu_instruction_master_granted_pcp_cpu_jtag_debug_module,
      pcp_cpu_instruction_master_qualified_request_pcp_cpu_jtag_debug_module => pcp_cpu_instruction_master_qualified_request_pcp_cpu_jtag_debug_module,
      pcp_cpu_instruction_master_read_data_valid_pcp_cpu_jtag_debug_module => pcp_cpu_instruction_master_read_data_valid_pcp_cpu_jtag_debug_module,
      pcp_cpu_instruction_master_requests_pcp_cpu_jtag_debug_module => pcp_cpu_instruction_master_requests_pcp_cpu_jtag_debug_module,
      pcp_cpu_jtag_debug_module_address => pcp_cpu_jtag_debug_module_address,
      pcp_cpu_jtag_debug_module_begintransfer => pcp_cpu_jtag_debug_module_begintransfer,
      pcp_cpu_jtag_debug_module_byteenable => pcp_cpu_jtag_debug_module_byteenable,
      pcp_cpu_jtag_debug_module_chipselect => pcp_cpu_jtag_debug_module_chipselect,
      pcp_cpu_jtag_debug_module_debugaccess => pcp_cpu_jtag_debug_module_debugaccess,
      pcp_cpu_jtag_debug_module_readdata_from_sa => pcp_cpu_jtag_debug_module_readdata_from_sa,
      pcp_cpu_jtag_debug_module_reset_n => pcp_cpu_jtag_debug_module_reset_n,
      pcp_cpu_jtag_debug_module_resetrequest_from_sa => pcp_cpu_jtag_debug_module_resetrequest_from_sa,
      pcp_cpu_jtag_debug_module_write => pcp_cpu_jtag_debug_module_write,
      pcp_cpu_jtag_debug_module_writedata => pcp_cpu_jtag_debug_module_writedata,
      clk => internal_clk90Meg,
      pcp_cpu_data_master_address_to_slave => pcp_cpu_data_master_address_to_slave,
      pcp_cpu_data_master_byteenable => pcp_cpu_data_master_byteenable,
      pcp_cpu_data_master_debugaccess => pcp_cpu_data_master_debugaccess,
      pcp_cpu_data_master_read => pcp_cpu_data_master_read,
      pcp_cpu_data_master_waitrequest => pcp_cpu_data_master_waitrequest,
      pcp_cpu_data_master_write => pcp_cpu_data_master_write,
      pcp_cpu_data_master_writedata => pcp_cpu_data_master_writedata,
      pcp_cpu_instruction_master_address_to_slave => pcp_cpu_instruction_master_address_to_slave,
      pcp_cpu_instruction_master_latency_counter => pcp_cpu_instruction_master_latency_counter,
      pcp_cpu_instruction_master_read => pcp_cpu_instruction_master_read,
      pcp_cpu_jtag_debug_module_readdata => pcp_cpu_jtag_debug_module_readdata,
      pcp_cpu_jtag_debug_module_resetrequest => pcp_cpu_jtag_debug_module_resetrequest,
      reset_n => clk90Meg_reset_n
    );


  --the_pcp_cpu_data_master, which is an e_instance
  the_pcp_cpu_data_master : pcp_cpu_data_master_arbitrator
    port map(
      pcp_cpu_data_master_address_to_slave => pcp_cpu_data_master_address_to_slave,
      pcp_cpu_data_master_dbs_address => pcp_cpu_data_master_dbs_address,
      pcp_cpu_data_master_dbs_write_16 => pcp_cpu_data_master_dbs_write_16,
      pcp_cpu_data_master_irq => pcp_cpu_data_master_irq,
      pcp_cpu_data_master_no_byte_enables_and_last_term => pcp_cpu_data_master_no_byte_enables_and_last_term,
      pcp_cpu_data_master_readdata => pcp_cpu_data_master_readdata,
      pcp_cpu_data_master_waitrequest => pcp_cpu_data_master_waitrequest,
      DBC3C40_SRAM_0_avalon_tristate_slave_wait_counter_eq_0 => DBC3C40_SRAM_0_avalon_tristate_slave_wait_counter_eq_0,
      OpenMAC_0_CMP_irq_from_sa => OpenMAC_0_CMP_irq_from_sa,
      OpenMAC_0_REG_irq_from_sa => OpenMAC_0_REG_irq_from_sa,
      OpenMAC_0_iBuf_readdata_from_sa => OpenMAC_0_iBuf_readdata_from_sa,
      OpenMAC_0_iBuf_wait_counter_eq_0 => OpenMAC_0_iBuf_wait_counter_eq_0,
      cfi_flash_0_s1_wait_counter_eq_0 => cfi_flash_0_s1_wait_counter_eq_0,
      cfi_flash_0_s1_wait_counter_eq_1 => cfi_flash_0_s1_wait_counter_eq_1,
      clk => internal_clk90Meg,
      clk90Meg => internal_clk90Meg,
      clk90Meg_reset_n => clk90Meg_reset_n,
      clock_crossing_0_s1_readdata_from_sa => clock_crossing_0_s1_readdata_from_sa,
      clock_crossing_0_s1_waitrequest_from_sa => clock_crossing_0_s1_waitrequest_from_sa,
      cnApi_Av2Av_0_pcp_readdata_from_sa => cnApi_Av2Av_0_pcp_readdata_from_sa,
      cnApi_Av2Av_0_pcp_wait_counter_eq_0 => cnApi_Av2Av_0_pcp_wait_counter_eq_0,
      d1_OpenMAC_0_iBuf_end_xfer => d1_OpenMAC_0_iBuf_end_xfer,
      d1_clock_crossing_0_s1_end_xfer => d1_clock_crossing_0_s1_end_xfer,
      d1_cnApi_Av2Av_0_pcp_end_xfer => d1_cnApi_Av2Av_0_pcp_end_xfer,
      d1_epcs_flash_controller_0_epcs_control_port_end_xfer => d1_epcs_flash_controller_0_epcs_control_port_end_xfer,
      d1_niosII_openMac_clock_0_in_end_xfer => d1_niosII_openMac_clock_0_in_end_xfer,
      d1_niosII_openMac_clock_1_in_end_xfer => d1_niosII_openMac_clock_1_in_end_xfer,
      d1_niosII_openMac_clock_2_in_end_xfer => d1_niosII_openMac_clock_2_in_end_xfer,
      d1_niosII_openMac_clock_3_in_end_xfer => d1_niosII_openMac_clock_3_in_end_xfer,
      d1_niosII_openMac_clock_4_in_end_xfer => d1_niosII_openMac_clock_4_in_end_xfer,
      d1_onchip_memory_0_s1_end_xfer => d1_onchip_memory_0_s1_end_xfer,
      d1_pcp_cpu_jtag_debug_module_end_xfer => d1_pcp_cpu_jtag_debug_module_end_xfer,
      d1_tri_state_bridge_0_avalon_slave_end_xfer => d1_tri_state_bridge_0_avalon_slave_end_xfer,
      epcs_flash_controller_0_epcs_control_port_irq_from_sa => epcs_flash_controller_0_epcs_control_port_irq_from_sa,
      epcs_flash_controller_0_epcs_control_port_readdata_from_sa => epcs_flash_controller_0_epcs_control_port_readdata_from_sa,
      incoming_tri_state_bridge_0_data => incoming_tri_state_bridge_0_data,
      incoming_tri_state_bridge_0_data_with_Xs_converted_to_0 => incoming_tri_state_bridge_0_data_with_Xs_converted_to_0,
      jtag_uart_0_avalon_jtag_slave_irq_from_sa => jtag_uart_0_avalon_jtag_slave_irq_from_sa,
      niosII_openMac_clock_0_in_readdata_from_sa => niosII_openMac_clock_0_in_readdata_from_sa,
      niosII_openMac_clock_0_in_waitrequest_from_sa => niosII_openMac_clock_0_in_waitrequest_from_sa,
      niosII_openMac_clock_1_in_readdata_from_sa => niosII_openMac_clock_1_in_readdata_from_sa,
      niosII_openMac_clock_1_in_waitrequest_from_sa => niosII_openMac_clock_1_in_waitrequest_from_sa,
      niosII_openMac_clock_2_in_readdata_from_sa => niosII_openMac_clock_2_in_readdata_from_sa,
      niosII_openMac_clock_2_in_waitrequest_from_sa => niosII_openMac_clock_2_in_waitrequest_from_sa,
      niosII_openMac_clock_3_in_readdata_from_sa => niosII_openMac_clock_3_in_readdata_from_sa,
      niosII_openMac_clock_3_in_waitrequest_from_sa => niosII_openMac_clock_3_in_waitrequest_from_sa,
      niosII_openMac_clock_4_in_readdata_from_sa => niosII_openMac_clock_4_in_readdata_from_sa,
      niosII_openMac_clock_4_in_waitrequest_from_sa => niosII_openMac_clock_4_in_waitrequest_from_sa,
      onchip_memory_0_s1_readdata_from_sa => onchip_memory_0_s1_readdata_from_sa,
      pcp_cpu_data_master_address => pcp_cpu_data_master_address,
      pcp_cpu_data_master_byteenable_DBC3C40_SRAM_0_avalon_tristate_slave => pcp_cpu_data_master_byteenable_DBC3C40_SRAM_0_avalon_tristate_slave,
      pcp_cpu_data_master_byteenable_cfi_flash_0_s1 => pcp_cpu_data_master_byteenable_cfi_flash_0_s1,
      pcp_cpu_data_master_byteenable_niosII_openMac_clock_2_in => pcp_cpu_data_master_byteenable_niosII_openMac_clock_2_in,
      pcp_cpu_data_master_granted_DBC3C40_SRAM_0_avalon_tristate_slave => pcp_cpu_data_master_granted_DBC3C40_SRAM_0_avalon_tristate_slave,
      pcp_cpu_data_master_granted_OpenMAC_0_iBuf => pcp_cpu_data_master_granted_OpenMAC_0_iBuf,
      pcp_cpu_data_master_granted_cfi_flash_0_s1 => pcp_cpu_data_master_granted_cfi_flash_0_s1,
      pcp_cpu_data_master_granted_clock_crossing_0_s1 => pcp_cpu_data_master_granted_clock_crossing_0_s1,
      pcp_cpu_data_master_granted_cnApi_Av2Av_0_pcp => pcp_cpu_data_master_granted_cnApi_Av2Av_0_pcp,
      pcp_cpu_data_master_granted_epcs_flash_controller_0_epcs_control_port => pcp_cpu_data_master_granted_epcs_flash_controller_0_epcs_control_port,
      pcp_cpu_data_master_granted_niosII_openMac_clock_0_in => pcp_cpu_data_master_granted_niosII_openMac_clock_0_in,
      pcp_cpu_data_master_granted_niosII_openMac_clock_1_in => pcp_cpu_data_master_granted_niosII_openMac_clock_1_in,
      pcp_cpu_data_master_granted_niosII_openMac_clock_2_in => pcp_cpu_data_master_granted_niosII_openMac_clock_2_in,
      pcp_cpu_data_master_granted_niosII_openMac_clock_3_in => pcp_cpu_data_master_granted_niosII_openMac_clock_3_in,
      pcp_cpu_data_master_granted_niosII_openMac_clock_4_in => pcp_cpu_data_master_granted_niosII_openMac_clock_4_in,
      pcp_cpu_data_master_granted_onchip_memory_0_s1 => pcp_cpu_data_master_granted_onchip_memory_0_s1,
      pcp_cpu_data_master_granted_pcp_cpu_jtag_debug_module => pcp_cpu_data_master_granted_pcp_cpu_jtag_debug_module,
      pcp_cpu_data_master_qualified_request_DBC3C40_SRAM_0_avalon_tristate_slave => pcp_cpu_data_master_qualified_request_DBC3C40_SRAM_0_avalon_tristate_slave,
      pcp_cpu_data_master_qualified_request_OpenMAC_0_iBuf => pcp_cpu_data_master_qualified_request_OpenMAC_0_iBuf,
      pcp_cpu_data_master_qualified_request_cfi_flash_0_s1 => pcp_cpu_data_master_qualified_request_cfi_flash_0_s1,
      pcp_cpu_data_master_qualified_request_clock_crossing_0_s1 => pcp_cpu_data_master_qualified_request_clock_crossing_0_s1,
      pcp_cpu_data_master_qualified_request_cnApi_Av2Av_0_pcp => pcp_cpu_data_master_qualified_request_cnApi_Av2Av_0_pcp,
      pcp_cpu_data_master_qualified_request_epcs_flash_controller_0_epcs_control_port => pcp_cpu_data_master_qualified_request_epcs_flash_controller_0_epcs_control_port,
      pcp_cpu_data_master_qualified_request_niosII_openMac_clock_0_in => pcp_cpu_data_master_qualified_request_niosII_openMac_clock_0_in,
      pcp_cpu_data_master_qualified_request_niosII_openMac_clock_1_in => pcp_cpu_data_master_qualified_request_niosII_openMac_clock_1_in,
      pcp_cpu_data_master_qualified_request_niosII_openMac_clock_2_in => pcp_cpu_data_master_qualified_request_niosII_openMac_clock_2_in,
      pcp_cpu_data_master_qualified_request_niosII_openMac_clock_3_in => pcp_cpu_data_master_qualified_request_niosII_openMac_clock_3_in,
      pcp_cpu_data_master_qualified_request_niosII_openMac_clock_4_in => pcp_cpu_data_master_qualified_request_niosII_openMac_clock_4_in,
      pcp_cpu_data_master_qualified_request_onchip_memory_0_s1 => pcp_cpu_data_master_qualified_request_onchip_memory_0_s1,
      pcp_cpu_data_master_qualified_request_pcp_cpu_jtag_debug_module => pcp_cpu_data_master_qualified_request_pcp_cpu_jtag_debug_module,
      pcp_cpu_data_master_read => pcp_cpu_data_master_read,
      pcp_cpu_data_master_read_data_valid_DBC3C40_SRAM_0_avalon_tristate_slave => pcp_cpu_data_master_read_data_valid_DBC3C40_SRAM_0_avalon_tristate_slave,
      pcp_cpu_data_master_read_data_valid_OpenMAC_0_iBuf => pcp_cpu_data_master_read_data_valid_OpenMAC_0_iBuf,
      pcp_cpu_data_master_read_data_valid_cfi_flash_0_s1 => pcp_cpu_data_master_read_data_valid_cfi_flash_0_s1,
      pcp_cpu_data_master_read_data_valid_clock_crossing_0_s1 => pcp_cpu_data_master_read_data_valid_clock_crossing_0_s1,
      pcp_cpu_data_master_read_data_valid_clock_crossing_0_s1_shift_register => pcp_cpu_data_master_read_data_valid_clock_crossing_0_s1_shift_register,
      pcp_cpu_data_master_read_data_valid_cnApi_Av2Av_0_pcp => pcp_cpu_data_master_read_data_valid_cnApi_Av2Av_0_pcp,
      pcp_cpu_data_master_read_data_valid_epcs_flash_controller_0_epcs_control_port => pcp_cpu_data_master_read_data_valid_epcs_flash_controller_0_epcs_control_port,
      pcp_cpu_data_master_read_data_valid_niosII_openMac_clock_0_in => pcp_cpu_data_master_read_data_valid_niosII_openMac_clock_0_in,
      pcp_cpu_data_master_read_data_valid_niosII_openMac_clock_1_in => pcp_cpu_data_master_read_data_valid_niosII_openMac_clock_1_in,
      pcp_cpu_data_master_read_data_valid_niosII_openMac_clock_2_in => pcp_cpu_data_master_read_data_valid_niosII_openMac_clock_2_in,
      pcp_cpu_data_master_read_data_valid_niosII_openMac_clock_3_in => pcp_cpu_data_master_read_data_valid_niosII_openMac_clock_3_in,
      pcp_cpu_data_master_read_data_valid_niosII_openMac_clock_4_in => pcp_cpu_data_master_read_data_valid_niosII_openMac_clock_4_in,
      pcp_cpu_data_master_read_data_valid_onchip_memory_0_s1 => pcp_cpu_data_master_read_data_valid_onchip_memory_0_s1,
      pcp_cpu_data_master_read_data_valid_pcp_cpu_jtag_debug_module => pcp_cpu_data_master_read_data_valid_pcp_cpu_jtag_debug_module,
      pcp_cpu_data_master_requests_DBC3C40_SRAM_0_avalon_tristate_slave => pcp_cpu_data_master_requests_DBC3C40_SRAM_0_avalon_tristate_slave,
      pcp_cpu_data_master_requests_OpenMAC_0_iBuf => pcp_cpu_data_master_requests_OpenMAC_0_iBuf,
      pcp_cpu_data_master_requests_cfi_flash_0_s1 => pcp_cpu_data_master_requests_cfi_flash_0_s1,
      pcp_cpu_data_master_requests_clock_crossing_0_s1 => pcp_cpu_data_master_requests_clock_crossing_0_s1,
      pcp_cpu_data_master_requests_cnApi_Av2Av_0_pcp => pcp_cpu_data_master_requests_cnApi_Av2Av_0_pcp,
      pcp_cpu_data_master_requests_epcs_flash_controller_0_epcs_control_port => pcp_cpu_data_master_requests_epcs_flash_controller_0_epcs_control_port,
      pcp_cpu_data_master_requests_niosII_openMac_clock_0_in => pcp_cpu_data_master_requests_niosII_openMac_clock_0_in,
      pcp_cpu_data_master_requests_niosII_openMac_clock_1_in => pcp_cpu_data_master_requests_niosII_openMac_clock_1_in,
      pcp_cpu_data_master_requests_niosII_openMac_clock_2_in => pcp_cpu_data_master_requests_niosII_openMac_clock_2_in,
      pcp_cpu_data_master_requests_niosII_openMac_clock_3_in => pcp_cpu_data_master_requests_niosII_openMac_clock_3_in,
      pcp_cpu_data_master_requests_niosII_openMac_clock_4_in => pcp_cpu_data_master_requests_niosII_openMac_clock_4_in,
      pcp_cpu_data_master_requests_onchip_memory_0_s1 => pcp_cpu_data_master_requests_onchip_memory_0_s1,
      pcp_cpu_data_master_requests_pcp_cpu_jtag_debug_module => pcp_cpu_data_master_requests_pcp_cpu_jtag_debug_module,
      pcp_cpu_data_master_write => pcp_cpu_data_master_write,
      pcp_cpu_data_master_writedata => pcp_cpu_data_master_writedata,
      pcp_cpu_jtag_debug_module_readdata_from_sa => pcp_cpu_jtag_debug_module_readdata_from_sa,
      registered_pcp_cpu_data_master_read_data_valid_DBC3C40_SRAM_0_avalon_tristate_slave => registered_pcp_cpu_data_master_read_data_valid_DBC3C40_SRAM_0_avalon_tristate_slave,
      registered_pcp_cpu_data_master_read_data_valid_cfi_flash_0_s1 => registered_pcp_cpu_data_master_read_data_valid_cfi_flash_0_s1,
      registered_pcp_cpu_data_master_read_data_valid_onchip_memory_0_s1 => registered_pcp_cpu_data_master_read_data_valid_onchip_memory_0_s1,
      reset_n => clk90Meg_reset_n,
      system_timer_s1_irq_from_sa => system_timer_s1_irq_from_sa
    );


  --the_pcp_cpu_instruction_master, which is an e_instance
  the_pcp_cpu_instruction_master : pcp_cpu_instruction_master_arbitrator
    port map(
      pcp_cpu_instruction_master_address_to_slave => pcp_cpu_instruction_master_address_to_slave,
      pcp_cpu_instruction_master_dbs_address => pcp_cpu_instruction_master_dbs_address,
      pcp_cpu_instruction_master_latency_counter => pcp_cpu_instruction_master_latency_counter,
      pcp_cpu_instruction_master_readdata => pcp_cpu_instruction_master_readdata,
      pcp_cpu_instruction_master_readdatavalid => pcp_cpu_instruction_master_readdatavalid,
      pcp_cpu_instruction_master_waitrequest => pcp_cpu_instruction_master_waitrequest,
      DBC3C40_SRAM_0_avalon_tristate_slave_wait_counter_eq_0 => DBC3C40_SRAM_0_avalon_tristate_slave_wait_counter_eq_0,
      cfi_flash_0_s1_wait_counter_eq_0 => cfi_flash_0_s1_wait_counter_eq_0,
      cfi_flash_0_s1_wait_counter_eq_1 => cfi_flash_0_s1_wait_counter_eq_1,
      clk => internal_clk90Meg,
      d1_epcs_flash_controller_0_epcs_control_port_end_xfer => d1_epcs_flash_controller_0_epcs_control_port_end_xfer,
      d1_onchip_memory_0_s1_end_xfer => d1_onchip_memory_0_s1_end_xfer,
      d1_pcp_cpu_jtag_debug_module_end_xfer => d1_pcp_cpu_jtag_debug_module_end_xfer,
      d1_tri_state_bridge_0_avalon_slave_end_xfer => d1_tri_state_bridge_0_avalon_slave_end_xfer,
      epcs_flash_controller_0_epcs_control_port_readdata_from_sa => epcs_flash_controller_0_epcs_control_port_readdata_from_sa,
      incoming_tri_state_bridge_0_data => incoming_tri_state_bridge_0_data,
      onchip_memory_0_s1_readdata_from_sa => onchip_memory_0_s1_readdata_from_sa,
      pcp_cpu_instruction_master_address => pcp_cpu_instruction_master_address,
      pcp_cpu_instruction_master_granted_DBC3C40_SRAM_0_avalon_tristate_slave => pcp_cpu_instruction_master_granted_DBC3C40_SRAM_0_avalon_tristate_slave,
      pcp_cpu_instruction_master_granted_cfi_flash_0_s1 => pcp_cpu_instruction_master_granted_cfi_flash_0_s1,
      pcp_cpu_instruction_master_granted_epcs_flash_controller_0_epcs_control_port => pcp_cpu_instruction_master_granted_epcs_flash_controller_0_epcs_control_port,
      pcp_cpu_instruction_master_granted_onchip_memory_0_s1 => pcp_cpu_instruction_master_granted_onchip_memory_0_s1,
      pcp_cpu_instruction_master_granted_pcp_cpu_jtag_debug_module => pcp_cpu_instruction_master_granted_pcp_cpu_jtag_debug_module,
      pcp_cpu_instruction_master_qualified_request_DBC3C40_SRAM_0_avalon_tristate_slave => pcp_cpu_instruction_master_qualified_request_DBC3C40_SRAM_0_avalon_tristate_slave,
      pcp_cpu_instruction_master_qualified_request_cfi_flash_0_s1 => pcp_cpu_instruction_master_qualified_request_cfi_flash_0_s1,
      pcp_cpu_instruction_master_qualified_request_epcs_flash_controller_0_epcs_control_port => pcp_cpu_instruction_master_qualified_request_epcs_flash_controller_0_epcs_control_port,
      pcp_cpu_instruction_master_qualified_request_onchip_memory_0_s1 => pcp_cpu_instruction_master_qualified_request_onchip_memory_0_s1,
      pcp_cpu_instruction_master_qualified_request_pcp_cpu_jtag_debug_module => pcp_cpu_instruction_master_qualified_request_pcp_cpu_jtag_debug_module,
      pcp_cpu_instruction_master_read => pcp_cpu_instruction_master_read,
      pcp_cpu_instruction_master_read_data_valid_DBC3C40_SRAM_0_avalon_tristate_slave => pcp_cpu_instruction_master_read_data_valid_DBC3C40_SRAM_0_avalon_tristate_slave,
      pcp_cpu_instruction_master_read_data_valid_cfi_flash_0_s1 => pcp_cpu_instruction_master_read_data_valid_cfi_flash_0_s1,
      pcp_cpu_instruction_master_read_data_valid_epcs_flash_controller_0_epcs_control_port => pcp_cpu_instruction_master_read_data_valid_epcs_flash_controller_0_epcs_control_port,
      pcp_cpu_instruction_master_read_data_valid_onchip_memory_0_s1 => pcp_cpu_instruction_master_read_data_valid_onchip_memory_0_s1,
      pcp_cpu_instruction_master_read_data_valid_pcp_cpu_jtag_debug_module => pcp_cpu_instruction_master_read_data_valid_pcp_cpu_jtag_debug_module,
      pcp_cpu_instruction_master_requests_DBC3C40_SRAM_0_avalon_tristate_slave => pcp_cpu_instruction_master_requests_DBC3C40_SRAM_0_avalon_tristate_slave,
      pcp_cpu_instruction_master_requests_cfi_flash_0_s1 => pcp_cpu_instruction_master_requests_cfi_flash_0_s1,
      pcp_cpu_instruction_master_requests_epcs_flash_controller_0_epcs_control_port => pcp_cpu_instruction_master_requests_epcs_flash_controller_0_epcs_control_port,
      pcp_cpu_instruction_master_requests_onchip_memory_0_s1 => pcp_cpu_instruction_master_requests_onchip_memory_0_s1,
      pcp_cpu_instruction_master_requests_pcp_cpu_jtag_debug_module => pcp_cpu_instruction_master_requests_pcp_cpu_jtag_debug_module,
      pcp_cpu_jtag_debug_module_readdata_from_sa => pcp_cpu_jtag_debug_module_readdata_from_sa,
      reset_n => clk90Meg_reset_n
    );


  --the_pcp_cpu, which is an e_ptf_instance
  the_pcp_cpu : pcp_cpu
    port map(
      d_address => pcp_cpu_data_master_address,
      d_byteenable => pcp_cpu_data_master_byteenable,
      d_read => pcp_cpu_data_master_read,
      d_write => pcp_cpu_data_master_write,
      d_writedata => pcp_cpu_data_master_writedata,
      i_address => pcp_cpu_instruction_master_address,
      i_read => pcp_cpu_instruction_master_read,
      jtag_debug_module_debugaccess_to_roms => pcp_cpu_data_master_debugaccess,
      jtag_debug_module_readdata => pcp_cpu_jtag_debug_module_readdata,
      jtag_debug_module_resetrequest => pcp_cpu_jtag_debug_module_resetrequest,
      clk => internal_clk90Meg,
      d_irq => pcp_cpu_data_master_irq,
      d_readdata => pcp_cpu_data_master_readdata,
      d_waitrequest => pcp_cpu_data_master_waitrequest,
      i_readdata => pcp_cpu_instruction_master_readdata,
      i_readdatavalid => pcp_cpu_instruction_master_readdatavalid,
      i_waitrequest => pcp_cpu_instruction_master_waitrequest,
      jtag_debug_module_address => pcp_cpu_jtag_debug_module_address,
      jtag_debug_module_begintransfer => pcp_cpu_jtag_debug_module_begintransfer,
      jtag_debug_module_byteenable => pcp_cpu_jtag_debug_module_byteenable,
      jtag_debug_module_debugaccess => pcp_cpu_jtag_debug_module_debugaccess,
      jtag_debug_module_select => pcp_cpu_jtag_debug_module_chipselect,
      jtag_debug_module_write => pcp_cpu_jtag_debug_module_write,
      jtag_debug_module_writedata => pcp_cpu_jtag_debug_module_writedata,
      reset_n => pcp_cpu_jtag_debug_module_reset_n
    );


  --the_portconf_pio_s1, which is an e_instance
  the_portconf_pio_s1 : portconf_pio_s1_arbitrator
    port map(
      clock_crossing_1_m1_granted_portconf_pio_s1 => clock_crossing_1_m1_granted_portconf_pio_s1,
      clock_crossing_1_m1_qualified_request_portconf_pio_s1 => clock_crossing_1_m1_qualified_request_portconf_pio_s1,
      clock_crossing_1_m1_read_data_valid_portconf_pio_s1 => clock_crossing_1_m1_read_data_valid_portconf_pio_s1,
      clock_crossing_1_m1_requests_portconf_pio_s1 => clock_crossing_1_m1_requests_portconf_pio_s1,
      d1_portconf_pio_s1_end_xfer => d1_portconf_pio_s1_end_xfer,
      portconf_pio_s1_address => portconf_pio_s1_address,
      portconf_pio_s1_chipselect => portconf_pio_s1_chipselect,
      portconf_pio_s1_readdata_from_sa => portconf_pio_s1_readdata_from_sa,
      portconf_pio_s1_reset_n => portconf_pio_s1_reset_n,
      portconf_pio_s1_write_n => portconf_pio_s1_write_n,
      portconf_pio_s1_writedata => portconf_pio_s1_writedata,
      clk => internal_clk50Meg,
      clock_crossing_1_m1_address_to_slave => clock_crossing_1_m1_address_to_slave,
      clock_crossing_1_m1_latency_counter => clock_crossing_1_m1_latency_counter,
      clock_crossing_1_m1_nativeaddress => clock_crossing_1_m1_nativeaddress,
      clock_crossing_1_m1_read => clock_crossing_1_m1_read,
      clock_crossing_1_m1_write => clock_crossing_1_m1_write,
      clock_crossing_1_m1_writedata => clock_crossing_1_m1_writedata,
      portconf_pio_s1_readdata => portconf_pio_s1_readdata,
      reset_n => clk50Meg_reset_n
    );


  --the_portconf_pio, which is an e_ptf_instance
  the_portconf_pio : portconf_pio
    port map(
      out_port => internal_out_port_from_the_portconf_pio,
      readdata => portconf_pio_s1_readdata,
      address => portconf_pio_s1_address,
      chipselect => portconf_pio_s1_chipselect,
      clk => internal_clk50Meg,
      in_port => in_port_to_the_portconf_pio,
      reset_n => portconf_pio_s1_reset_n,
      write_n => portconf_pio_s1_write_n,
      writedata => portconf_pio_s1_writedata
    );


  --the_remote_update_cycloneiii_0_s1, which is an e_instance
  the_remote_update_cycloneiii_0_s1 : remote_update_cycloneiii_0_s1_arbitrator
    port map(
      d1_remote_update_cycloneiii_0_s1_end_xfer => d1_remote_update_cycloneiii_0_s1_end_xfer,
      niosII_openMac_clock_4_out_granted_remote_update_cycloneiii_0_s1 => niosII_openMac_clock_4_out_granted_remote_update_cycloneiii_0_s1,
      niosII_openMac_clock_4_out_qualified_request_remote_update_cycloneiii_0_s1 => niosII_openMac_clock_4_out_qualified_request_remote_update_cycloneiii_0_s1,
      niosII_openMac_clock_4_out_read_data_valid_remote_update_cycloneiii_0_s1 => niosII_openMac_clock_4_out_read_data_valid_remote_update_cycloneiii_0_s1,
      niosII_openMac_clock_4_out_requests_remote_update_cycloneiii_0_s1 => niosII_openMac_clock_4_out_requests_remote_update_cycloneiii_0_s1,
      remote_update_cycloneiii_0_s1_address => remote_update_cycloneiii_0_s1_address,
      remote_update_cycloneiii_0_s1_chipselect => remote_update_cycloneiii_0_s1_chipselect,
      remote_update_cycloneiii_0_s1_read => remote_update_cycloneiii_0_s1_read,
      remote_update_cycloneiii_0_s1_readdata_from_sa => remote_update_cycloneiii_0_s1_readdata_from_sa,
      remote_update_cycloneiii_0_s1_reset => remote_update_cycloneiii_0_s1_reset,
      remote_update_cycloneiii_0_s1_waitrequest_from_sa => remote_update_cycloneiii_0_s1_waitrequest_from_sa,
      remote_update_cycloneiii_0_s1_write => remote_update_cycloneiii_0_s1_write,
      remote_update_cycloneiii_0_s1_writedata => remote_update_cycloneiii_0_s1_writedata,
      clk => internal_clk25Meg,
      niosII_openMac_clock_4_out_address_to_slave => niosII_openMac_clock_4_out_address_to_slave,
      niosII_openMac_clock_4_out_nativeaddress => niosII_openMac_clock_4_out_nativeaddress,
      niosII_openMac_clock_4_out_read => niosII_openMac_clock_4_out_read,
      niosII_openMac_clock_4_out_write => niosII_openMac_clock_4_out_write,
      niosII_openMac_clock_4_out_writedata => niosII_openMac_clock_4_out_writedata,
      remote_update_cycloneiii_0_s1_readdata => remote_update_cycloneiii_0_s1_readdata,
      remote_update_cycloneiii_0_s1_waitrequest => remote_update_cycloneiii_0_s1_waitrequest,
      reset_n => clk25Meg_reset_n
    );


  --the_remote_update_cycloneiii_0, which is an e_ptf_instance
  the_remote_update_cycloneiii_0 : remote_update_cycloneiii_0
    port map(
      readdata => remote_update_cycloneiii_0_s1_readdata,
      waitrequest => remote_update_cycloneiii_0_s1_waitrequest,
      address => remote_update_cycloneiii_0_s1_address,
      chipselect => remote_update_cycloneiii_0_s1_chipselect,
      clk => internal_clk25Meg,
      read => remote_update_cycloneiii_0_s1_read,
      reset => remote_update_cycloneiii_0_s1_reset,
      write => remote_update_cycloneiii_0_s1_write,
      writedata => remote_update_cycloneiii_0_s1_writedata
    );


  --the_sdram_0_s1, which is an e_instance
  the_sdram_0_s1 : sdram_0_s1_arbitrator
    port map(
      ap_cpu_data_master_granted_sdram_0_s1 => ap_cpu_data_master_granted_sdram_0_s1,
      ap_cpu_data_master_qualified_request_sdram_0_s1 => ap_cpu_data_master_qualified_request_sdram_0_s1,
      ap_cpu_data_master_read_data_valid_sdram_0_s1 => ap_cpu_data_master_read_data_valid_sdram_0_s1,
      ap_cpu_data_master_read_data_valid_sdram_0_s1_shift_register => ap_cpu_data_master_read_data_valid_sdram_0_s1_shift_register,
      ap_cpu_data_master_requests_sdram_0_s1 => ap_cpu_data_master_requests_sdram_0_s1,
      ap_cpu_instruction_master_granted_sdram_0_s1 => ap_cpu_instruction_master_granted_sdram_0_s1,
      ap_cpu_instruction_master_qualified_request_sdram_0_s1 => ap_cpu_instruction_master_qualified_request_sdram_0_s1,
      ap_cpu_instruction_master_read_data_valid_sdram_0_s1 => ap_cpu_instruction_master_read_data_valid_sdram_0_s1,
      ap_cpu_instruction_master_read_data_valid_sdram_0_s1_shift_register => ap_cpu_instruction_master_read_data_valid_sdram_0_s1_shift_register,
      ap_cpu_instruction_master_requests_sdram_0_s1 => ap_cpu_instruction_master_requests_sdram_0_s1,
      d1_sdram_0_s1_end_xfer => d1_sdram_0_s1_end_xfer,
      sdram_0_s1_address => sdram_0_s1_address,
      sdram_0_s1_byteenable_n => sdram_0_s1_byteenable_n,
      sdram_0_s1_chipselect => sdram_0_s1_chipselect,
      sdram_0_s1_read_n => sdram_0_s1_read_n,
      sdram_0_s1_readdata_from_sa => sdram_0_s1_readdata_from_sa,
      sdram_0_s1_reset_n => sdram_0_s1_reset_n,
      sdram_0_s1_waitrequest_from_sa => sdram_0_s1_waitrequest_from_sa,
      sdram_0_s1_write_n => sdram_0_s1_write_n,
      sdram_0_s1_writedata => sdram_0_s1_writedata,
      ap_cpu_data_master_address_to_slave => ap_cpu_data_master_address_to_slave,
      ap_cpu_data_master_byteenable => ap_cpu_data_master_byteenable,
      ap_cpu_data_master_read => ap_cpu_data_master_read,
      ap_cpu_data_master_waitrequest => ap_cpu_data_master_waitrequest,
      ap_cpu_data_master_write => ap_cpu_data_master_write,
      ap_cpu_data_master_writedata => ap_cpu_data_master_writedata,
      ap_cpu_instruction_master_address_to_slave => ap_cpu_instruction_master_address_to_slave,
      ap_cpu_instruction_master_latency_counter => ap_cpu_instruction_master_latency_counter,
      ap_cpu_instruction_master_read => ap_cpu_instruction_master_read,
      clk => internal_clk90Meg,
      reset_n => clk90Meg_reset_n,
      sdram_0_s1_readdata => sdram_0_s1_readdata,
      sdram_0_s1_readdatavalid => sdram_0_s1_readdatavalid,
      sdram_0_s1_waitrequest => sdram_0_s1_waitrequest
    );


  --the_sdram_0, which is an e_ptf_instance
  the_sdram_0 : sdram_0
    port map(
      za_data => sdram_0_s1_readdata,
      za_valid => sdram_0_s1_readdatavalid,
      za_waitrequest => sdram_0_s1_waitrequest,
      zs_addr => internal_zs_addr_from_the_sdram_0,
      zs_ba => internal_zs_ba_from_the_sdram_0,
      zs_cas_n => internal_zs_cas_n_from_the_sdram_0,
      zs_cke => internal_zs_cke_from_the_sdram_0,
      zs_cs_n => internal_zs_cs_n_from_the_sdram_0,
      zs_dq => zs_dq_to_and_from_the_sdram_0,
      zs_dqm => internal_zs_dqm_from_the_sdram_0,
      zs_ras_n => internal_zs_ras_n_from_the_sdram_0,
      zs_we_n => internal_zs_we_n_from_the_sdram_0,
      az_addr => sdram_0_s1_address,
      az_be_n => sdram_0_s1_byteenable_n,
      az_cs => sdram_0_s1_chipselect,
      az_data => sdram_0_s1_writedata,
      az_rd_n => sdram_0_s1_read_n,
      az_wr_n => sdram_0_s1_write_n,
      clk => internal_clk90Meg,
      reset_n => sdram_0_s1_reset_n
    );


  --the_status_led_pio_s1, which is an e_instance
  the_status_led_pio_s1 : status_led_pio_s1_arbitrator
    port map(
      clock_crossing_0_m1_granted_status_led_pio_s1 => clock_crossing_0_m1_granted_status_led_pio_s1,
      clock_crossing_0_m1_qualified_request_status_led_pio_s1 => clock_crossing_0_m1_qualified_request_status_led_pio_s1,
      clock_crossing_0_m1_read_data_valid_status_led_pio_s1 => clock_crossing_0_m1_read_data_valid_status_led_pio_s1,
      clock_crossing_0_m1_requests_status_led_pio_s1 => clock_crossing_0_m1_requests_status_led_pio_s1,
      d1_status_led_pio_s1_end_xfer => d1_status_led_pio_s1_end_xfer,
      status_led_pio_s1_address => status_led_pio_s1_address,
      status_led_pio_s1_chipselect => status_led_pio_s1_chipselect,
      status_led_pio_s1_readdata_from_sa => status_led_pio_s1_readdata_from_sa,
      status_led_pio_s1_reset_n => status_led_pio_s1_reset_n,
      status_led_pio_s1_write_n => status_led_pio_s1_write_n,
      status_led_pio_s1_writedata => status_led_pio_s1_writedata,
      clk => internal_clk50Meg,
      clock_crossing_0_m1_address_to_slave => clock_crossing_0_m1_address_to_slave,
      clock_crossing_0_m1_byteenable => clock_crossing_0_m1_byteenable,
      clock_crossing_0_m1_latency_counter => clock_crossing_0_m1_latency_counter,
      clock_crossing_0_m1_nativeaddress => clock_crossing_0_m1_nativeaddress,
      clock_crossing_0_m1_read => clock_crossing_0_m1_read,
      clock_crossing_0_m1_write => clock_crossing_0_m1_write,
      clock_crossing_0_m1_writedata => clock_crossing_0_m1_writedata,
      reset_n => clk50Meg_reset_n,
      status_led_pio_s1_readdata => status_led_pio_s1_readdata
    );


  --the_status_led_pio, which is an e_ptf_instance
  the_status_led_pio : status_led_pio
    port map(
      out_port => internal_out_port_from_the_status_led_pio,
      readdata => status_led_pio_s1_readdata,
      address => status_led_pio_s1_address,
      chipselect => status_led_pio_s1_chipselect,
      clk => internal_clk50Meg,
      reset_n => status_led_pio_s1_reset_n,
      write_n => status_led_pio_s1_write_n,
      writedata => status_led_pio_s1_writedata
    );


  --the_sync_irq_s1, which is an e_instance
  the_sync_irq_s1 : sync_irq_s1_arbitrator
    port map(
      clock_crossing_1_m1_granted_sync_irq_s1 => clock_crossing_1_m1_granted_sync_irq_s1,
      clock_crossing_1_m1_qualified_request_sync_irq_s1 => clock_crossing_1_m1_qualified_request_sync_irq_s1,
      clock_crossing_1_m1_read_data_valid_sync_irq_s1 => clock_crossing_1_m1_read_data_valid_sync_irq_s1,
      clock_crossing_1_m1_requests_sync_irq_s1 => clock_crossing_1_m1_requests_sync_irq_s1,
      d1_sync_irq_s1_end_xfer => d1_sync_irq_s1_end_xfer,
      sync_irq_s1_address => sync_irq_s1_address,
      sync_irq_s1_chipselect => sync_irq_s1_chipselect,
      sync_irq_s1_irq_from_sa => sync_irq_s1_irq_from_sa,
      sync_irq_s1_readdata_from_sa => sync_irq_s1_readdata_from_sa,
      sync_irq_s1_reset_n => sync_irq_s1_reset_n,
      sync_irq_s1_write_n => sync_irq_s1_write_n,
      sync_irq_s1_writedata => sync_irq_s1_writedata,
      clk => internal_clk50Meg,
      clock_crossing_1_m1_address_to_slave => clock_crossing_1_m1_address_to_slave,
      clock_crossing_1_m1_latency_counter => clock_crossing_1_m1_latency_counter,
      clock_crossing_1_m1_nativeaddress => clock_crossing_1_m1_nativeaddress,
      clock_crossing_1_m1_read => clock_crossing_1_m1_read,
      clock_crossing_1_m1_write => clock_crossing_1_m1_write,
      clock_crossing_1_m1_writedata => clock_crossing_1_m1_writedata,
      reset_n => clk50Meg_reset_n,
      sync_irq_s1_irq => sync_irq_s1_irq,
      sync_irq_s1_readdata => sync_irq_s1_readdata
    );


  --the_sync_irq, which is an e_ptf_instance
  the_sync_irq : sync_irq
    port map(
      irq => sync_irq_s1_irq,
      readdata => sync_irq_s1_readdata,
      address => sync_irq_s1_address,
      chipselect => sync_irq_s1_chipselect,
      clk => internal_clk50Meg,
      in_port => in_port_to_the_sync_irq,
      reset_n => sync_irq_s1_reset_n,
      write_n => sync_irq_s1_write_n,
      writedata => sync_irq_s1_writedata
    );


  --the_sysid_control_slave, which is an e_instance
  the_sysid_control_slave : sysid_control_slave_arbitrator
    port map(
      clock_crossing_0_m1_granted_sysid_control_slave => clock_crossing_0_m1_granted_sysid_control_slave,
      clock_crossing_0_m1_qualified_request_sysid_control_slave => clock_crossing_0_m1_qualified_request_sysid_control_slave,
      clock_crossing_0_m1_read_data_valid_sysid_control_slave => clock_crossing_0_m1_read_data_valid_sysid_control_slave,
      clock_crossing_0_m1_requests_sysid_control_slave => clock_crossing_0_m1_requests_sysid_control_slave,
      clock_crossing_1_m1_granted_sysid_control_slave => clock_crossing_1_m1_granted_sysid_control_slave,
      clock_crossing_1_m1_qualified_request_sysid_control_slave => clock_crossing_1_m1_qualified_request_sysid_control_slave,
      clock_crossing_1_m1_read_data_valid_sysid_control_slave => clock_crossing_1_m1_read_data_valid_sysid_control_slave,
      clock_crossing_1_m1_requests_sysid_control_slave => clock_crossing_1_m1_requests_sysid_control_slave,
      d1_sysid_control_slave_end_xfer => d1_sysid_control_slave_end_xfer,
      sysid_control_slave_address => sysid_control_slave_address,
      sysid_control_slave_readdata_from_sa => sysid_control_slave_readdata_from_sa,
      clk => internal_clk50Meg,
      clock_crossing_0_m1_address_to_slave => clock_crossing_0_m1_address_to_slave,
      clock_crossing_0_m1_latency_counter => clock_crossing_0_m1_latency_counter,
      clock_crossing_0_m1_nativeaddress => clock_crossing_0_m1_nativeaddress,
      clock_crossing_0_m1_read => clock_crossing_0_m1_read,
      clock_crossing_0_m1_write => clock_crossing_0_m1_write,
      clock_crossing_1_m1_address_to_slave => clock_crossing_1_m1_address_to_slave,
      clock_crossing_1_m1_latency_counter => clock_crossing_1_m1_latency_counter,
      clock_crossing_1_m1_nativeaddress => clock_crossing_1_m1_nativeaddress,
      clock_crossing_1_m1_read => clock_crossing_1_m1_read,
      clock_crossing_1_m1_write => clock_crossing_1_m1_write,
      reset_n => clk50Meg_reset_n,
      sysid_control_slave_readdata => sysid_control_slave_readdata
    );


  --the_sysid, which is an e_ptf_instance
  the_sysid : sysid
    port map(
      readdata => sysid_control_slave_readdata,
      address => sysid_control_slave_address
    );


  --the_system_timer_s1, which is an e_instance
  the_system_timer_s1 : system_timer_s1_arbitrator
    port map(
      clock_crossing_0_m1_granted_system_timer_s1 => clock_crossing_0_m1_granted_system_timer_s1,
      clock_crossing_0_m1_qualified_request_system_timer_s1 => clock_crossing_0_m1_qualified_request_system_timer_s1,
      clock_crossing_0_m1_read_data_valid_system_timer_s1 => clock_crossing_0_m1_read_data_valid_system_timer_s1,
      clock_crossing_0_m1_requests_system_timer_s1 => clock_crossing_0_m1_requests_system_timer_s1,
      d1_system_timer_s1_end_xfer => d1_system_timer_s1_end_xfer,
      system_timer_s1_address => system_timer_s1_address,
      system_timer_s1_chipselect => system_timer_s1_chipselect,
      system_timer_s1_irq_from_sa => system_timer_s1_irq_from_sa,
      system_timer_s1_readdata_from_sa => system_timer_s1_readdata_from_sa,
      system_timer_s1_reset_n => system_timer_s1_reset_n,
      system_timer_s1_write_n => system_timer_s1_write_n,
      system_timer_s1_writedata => system_timer_s1_writedata,
      clk => internal_clk50Meg,
      clock_crossing_0_m1_address_to_slave => clock_crossing_0_m1_address_to_slave,
      clock_crossing_0_m1_latency_counter => clock_crossing_0_m1_latency_counter,
      clock_crossing_0_m1_nativeaddress => clock_crossing_0_m1_nativeaddress,
      clock_crossing_0_m1_read => clock_crossing_0_m1_read,
      clock_crossing_0_m1_write => clock_crossing_0_m1_write,
      clock_crossing_0_m1_writedata => clock_crossing_0_m1_writedata,
      reset_n => clk50Meg_reset_n,
      system_timer_s1_irq => system_timer_s1_irq,
      system_timer_s1_readdata => system_timer_s1_readdata
    );


  --the_system_timer, which is an e_ptf_instance
  the_system_timer : system_timer
    port map(
      irq => system_timer_s1_irq,
      readdata => system_timer_s1_readdata,
      address => system_timer_s1_address,
      chipselect => system_timer_s1_chipselect,
      clk => internal_clk50Meg,
      reset_n => system_timer_s1_reset_n,
      write_n => system_timer_s1_write_n,
      writedata => system_timer_s1_writedata
    );


  --the_system_timer_ap_s1, which is an e_instance
  the_system_timer_ap_s1 : system_timer_ap_s1_arbitrator
    port map(
      clock_crossing_1_m1_granted_system_timer_ap_s1 => clock_crossing_1_m1_granted_system_timer_ap_s1,
      clock_crossing_1_m1_qualified_request_system_timer_ap_s1 => clock_crossing_1_m1_qualified_request_system_timer_ap_s1,
      clock_crossing_1_m1_read_data_valid_system_timer_ap_s1 => clock_crossing_1_m1_read_data_valid_system_timer_ap_s1,
      clock_crossing_1_m1_requests_system_timer_ap_s1 => clock_crossing_1_m1_requests_system_timer_ap_s1,
      d1_system_timer_ap_s1_end_xfer => d1_system_timer_ap_s1_end_xfer,
      system_timer_ap_s1_address => system_timer_ap_s1_address,
      system_timer_ap_s1_chipselect => system_timer_ap_s1_chipselect,
      system_timer_ap_s1_irq_from_sa => system_timer_ap_s1_irq_from_sa,
      system_timer_ap_s1_readdata_from_sa => system_timer_ap_s1_readdata_from_sa,
      system_timer_ap_s1_reset_n => system_timer_ap_s1_reset_n,
      system_timer_ap_s1_write_n => system_timer_ap_s1_write_n,
      system_timer_ap_s1_writedata => system_timer_ap_s1_writedata,
      clk => internal_clk50Meg,
      clock_crossing_1_m1_address_to_slave => clock_crossing_1_m1_address_to_slave,
      clock_crossing_1_m1_latency_counter => clock_crossing_1_m1_latency_counter,
      clock_crossing_1_m1_nativeaddress => clock_crossing_1_m1_nativeaddress,
      clock_crossing_1_m1_read => clock_crossing_1_m1_read,
      clock_crossing_1_m1_write => clock_crossing_1_m1_write,
      clock_crossing_1_m1_writedata => clock_crossing_1_m1_writedata,
      reset_n => clk50Meg_reset_n,
      system_timer_ap_s1_irq => system_timer_ap_s1_irq,
      system_timer_ap_s1_readdata => system_timer_ap_s1_readdata
    );


  --the_system_timer_ap, which is an e_ptf_instance
  the_system_timer_ap : system_timer_ap
    port map(
      irq => system_timer_ap_s1_irq,
      readdata => system_timer_ap_s1_readdata,
      address => system_timer_ap_s1_address,
      chipselect => system_timer_ap_s1_chipselect,
      clk => internal_clk50Meg,
      reset_n => system_timer_ap_s1_reset_n,
      write_n => system_timer_ap_s1_write_n,
      writedata => system_timer_ap_s1_writedata
    );


  --the_tri_state_bridge_0_avalon_slave, which is an e_instance
  the_tri_state_bridge_0_avalon_slave : tri_state_bridge_0_avalon_slave_arbitrator
    port map(
      DBC3C40_SRAM_0_avalon_tristate_slave_wait_counter_eq_0 => DBC3C40_SRAM_0_avalon_tristate_slave_wait_counter_eq_0,
      ben_to_the_DBC3C40_SRAM_0 => internal_ben_to_the_DBC3C40_SRAM_0,
      cfi_flash_0_s1_wait_counter_eq_0 => cfi_flash_0_s1_wait_counter_eq_0,
      cfi_flash_0_s1_wait_counter_eq_1 => cfi_flash_0_s1_wait_counter_eq_1,
      d1_tri_state_bridge_0_avalon_slave_end_xfer => d1_tri_state_bridge_0_avalon_slave_end_xfer,
      incoming_tri_state_bridge_0_data => incoming_tri_state_bridge_0_data,
      incoming_tri_state_bridge_0_data_with_Xs_converted_to_0 => incoming_tri_state_bridge_0_data_with_Xs_converted_to_0,
      ncs_to_the_DBC3C40_SRAM_0 => internal_ncs_to_the_DBC3C40_SRAM_0,
      pcp_cpu_data_master_byteenable_DBC3C40_SRAM_0_avalon_tristate_slave => pcp_cpu_data_master_byteenable_DBC3C40_SRAM_0_avalon_tristate_slave,
      pcp_cpu_data_master_byteenable_cfi_flash_0_s1 => pcp_cpu_data_master_byteenable_cfi_flash_0_s1,
      pcp_cpu_data_master_granted_DBC3C40_SRAM_0_avalon_tristate_slave => pcp_cpu_data_master_granted_DBC3C40_SRAM_0_avalon_tristate_slave,
      pcp_cpu_data_master_granted_cfi_flash_0_s1 => pcp_cpu_data_master_granted_cfi_flash_0_s1,
      pcp_cpu_data_master_qualified_request_DBC3C40_SRAM_0_avalon_tristate_slave => pcp_cpu_data_master_qualified_request_DBC3C40_SRAM_0_avalon_tristate_slave,
      pcp_cpu_data_master_qualified_request_cfi_flash_0_s1 => pcp_cpu_data_master_qualified_request_cfi_flash_0_s1,
      pcp_cpu_data_master_read_data_valid_DBC3C40_SRAM_0_avalon_tristate_slave => pcp_cpu_data_master_read_data_valid_DBC3C40_SRAM_0_avalon_tristate_slave,
      pcp_cpu_data_master_read_data_valid_cfi_flash_0_s1 => pcp_cpu_data_master_read_data_valid_cfi_flash_0_s1,
      pcp_cpu_data_master_requests_DBC3C40_SRAM_0_avalon_tristate_slave => pcp_cpu_data_master_requests_DBC3C40_SRAM_0_avalon_tristate_slave,
      pcp_cpu_data_master_requests_cfi_flash_0_s1 => pcp_cpu_data_master_requests_cfi_flash_0_s1,
      pcp_cpu_instruction_master_granted_DBC3C40_SRAM_0_avalon_tristate_slave => pcp_cpu_instruction_master_granted_DBC3C40_SRAM_0_avalon_tristate_slave,
      pcp_cpu_instruction_master_granted_cfi_flash_0_s1 => pcp_cpu_instruction_master_granted_cfi_flash_0_s1,
      pcp_cpu_instruction_master_qualified_request_DBC3C40_SRAM_0_avalon_tristate_slave => pcp_cpu_instruction_master_qualified_request_DBC3C40_SRAM_0_avalon_tristate_slave,
      pcp_cpu_instruction_master_qualified_request_cfi_flash_0_s1 => pcp_cpu_instruction_master_qualified_request_cfi_flash_0_s1,
      pcp_cpu_instruction_master_read_data_valid_DBC3C40_SRAM_0_avalon_tristate_slave => pcp_cpu_instruction_master_read_data_valid_DBC3C40_SRAM_0_avalon_tristate_slave,
      pcp_cpu_instruction_master_read_data_valid_cfi_flash_0_s1 => pcp_cpu_instruction_master_read_data_valid_cfi_flash_0_s1,
      pcp_cpu_instruction_master_requests_DBC3C40_SRAM_0_avalon_tristate_slave => pcp_cpu_instruction_master_requests_DBC3C40_SRAM_0_avalon_tristate_slave,
      pcp_cpu_instruction_master_requests_cfi_flash_0_s1 => pcp_cpu_instruction_master_requests_cfi_flash_0_s1,
      registered_pcp_cpu_data_master_read_data_valid_DBC3C40_SRAM_0_avalon_tristate_slave => registered_pcp_cpu_data_master_read_data_valid_DBC3C40_SRAM_0_avalon_tristate_slave,
      registered_pcp_cpu_data_master_read_data_valid_cfi_flash_0_s1 => registered_pcp_cpu_data_master_read_data_valid_cfi_flash_0_s1,
      select_n_to_the_cfi_flash_0 => internal_select_n_to_the_cfi_flash_0,
      tri_state_bridge_0_address => internal_tri_state_bridge_0_address,
      tri_state_bridge_0_data => tri_state_bridge_0_data,
      tri_state_bridge_0_readn => internal_tri_state_bridge_0_readn,
      tri_state_bridge_0_writen => internal_tri_state_bridge_0_writen,
      clk => internal_clk90Meg,
      pcp_cpu_data_master_address_to_slave => pcp_cpu_data_master_address_to_slave,
      pcp_cpu_data_master_byteenable => pcp_cpu_data_master_byteenable,
      pcp_cpu_data_master_dbs_address => pcp_cpu_data_master_dbs_address,
      pcp_cpu_data_master_dbs_write_16 => pcp_cpu_data_master_dbs_write_16,
      pcp_cpu_data_master_no_byte_enables_and_last_term => pcp_cpu_data_master_no_byte_enables_and_last_term,
      pcp_cpu_data_master_read => pcp_cpu_data_master_read,
      pcp_cpu_data_master_write => pcp_cpu_data_master_write,
      pcp_cpu_instruction_master_address_to_slave => pcp_cpu_instruction_master_address_to_slave,
      pcp_cpu_instruction_master_dbs_address => pcp_cpu_instruction_master_dbs_address,
      pcp_cpu_instruction_master_latency_counter => pcp_cpu_instruction_master_latency_counter,
      pcp_cpu_instruction_master_read => pcp_cpu_instruction_master_read,
      reset_n => clk90Meg_reset_n
    );


  --reset is asserted asynchronously and deasserted synchronously
  niosII_openMac_reset_clk50Meg_domain_synch : niosII_openMac_reset_clk50Meg_domain_synch_module
    port map(
      data_out => clk50Meg_reset_n,
      clk => internal_clk50Meg,
      data_in => module_input12,
      reset_n => reset_n_sources
    );

  module_input12 <= std_logic'('1');

  --reset sources mux, which is an e_mux
  reset_n_sources <= Vector_To_Std_Logic(NOT ((((((((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT reset_n))) OR std_logic_vector'("00000000000000000000000000000000")) OR std_logic_vector'("00000000000000000000000000000000")) OR std_logic_vector'("00000000000000000000000000000000")) OR (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(ap_cpu_jtag_debug_module_resetrequest_from_sa)))) OR (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(ap_cpu_jtag_debug_module_resetrequest_from_sa)))) OR (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pcp_cpu_jtag_debug_module_resetrequest_from_sa)))) OR (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pcp_cpu_jtag_debug_module_resetrequest_from_sa)))) OR std_logic_vector'("00000000000000000000000000000000"))));
  --reset is asserted asynchronously and deasserted synchronously
  niosII_openMac_reset_clk90Meg_domain_synch : niosII_openMac_reset_clk90Meg_domain_synch_module
    port map(
      data_out => clk90Meg_reset_n,
      clk => internal_clk90Meg,
      data_in => module_input13,
      reset_n => reset_n_sources
    );

  module_input13 <= std_logic'('1');

  --reset is asserted asynchronously and deasserted synchronously
  niosII_openMac_reset_clk_0_domain_synch : niosII_openMac_reset_clk_0_domain_synch_module
    port map(
      data_out => clk_0_reset_n,
      clk => clk_0,
      data_in => module_input14,
      reset_n => reset_n_sources
    );

  module_input14 <= std_logic'('1');

  --reset is asserted asynchronously and deasserted synchronously
  niosII_openMac_reset_clk25Meg_domain_synch : niosII_openMac_reset_clk25Meg_domain_synch_module
    port map(
      data_out => clk25Meg_reset_n,
      clk => internal_clk25Meg,
      data_in => module_input15,
      reset_n => reset_n_sources
    );

  module_input15 <= std_logic'('1');

  --clock_crossing_0_m1_endofpacket of type endofpacket does not connect to anything so wire it to default (0)
  clock_crossing_0_m1_endofpacket <= std_logic'('0');
  --clock_crossing_1_m1_endofpacket of type endofpacket does not connect to anything so wire it to default (0)
  clock_crossing_1_m1_endofpacket <= std_logic'('0');
  --niosII_openMac_clock_0_out_endofpacket of type endofpacket does not connect to anything so wire it to default (0)
  niosII_openMac_clock_0_out_endofpacket <= std_logic'('0');
  --niosII_openMac_clock_1_out_endofpacket of type endofpacket does not connect to anything so wire it to default (0)
  niosII_openMac_clock_1_out_endofpacket <= std_logic'('0');
  --niosII_openMac_clock_2_out_endofpacket of type endofpacket does not connect to anything so wire it to default (0)
  niosII_openMac_clock_2_out_endofpacket <= std_logic'('0');
  --niosII_openMac_clock_3_out_endofpacket of type endofpacket does not connect to anything so wire it to default (0)
  niosII_openMac_clock_3_out_endofpacket <= std_logic'('0');
  --niosII_openMac_clock_4_out_endofpacket of type endofpacket does not connect to anything so wire it to default (0)
  niosII_openMac_clock_4_out_endofpacket <= std_logic'('0');
  --vhdl renameroo for output signals
  ben_to_the_DBC3C40_SRAM_0 <= internal_ben_to_the_DBC3C40_SRAM_0;
  --vhdl renameroo for output signals
  clk25Meg <= internal_clk25Meg;
  --vhdl renameroo for output signals
  clk50Meg <= internal_clk50Meg;
  --vhdl renameroo for output signals
  clk90Meg <= internal_clk90Meg;
  --vhdl renameroo for output signals
  dclk_from_the_epcs_flash_controller_0 <= internal_dclk_from_the_epcs_flash_controller_0;
  --vhdl renameroo for output signals
  locked_from_the_altpll_0 <= internal_locked_from_the_altpll_0;
  --vhdl renameroo for output signals
  mii_Clk_from_the_OpenMAC_0 <= internal_mii_Clk_from_the_OpenMAC_0;
  --vhdl renameroo for output signals
  mii_Do_from_the_OpenMAC_0 <= internal_mii_Do_from_the_OpenMAC_0;
  --vhdl renameroo for output signals
  mii_Doe_from_the_OpenMAC_0 <= internal_mii_Doe_from_the_OpenMAC_0;
  --vhdl renameroo for output signals
  mii_nResetOut_from_the_OpenMAC_0 <= internal_mii_nResetOut_from_the_OpenMAC_0;
  --vhdl renameroo for output signals
  ncs_to_the_DBC3C40_SRAM_0 <= internal_ncs_to_the_DBC3C40_SRAM_0;
  --vhdl renameroo for output signals
  out_port_from_the_irq_gen <= internal_out_port_from_the_irq_gen;
  --vhdl renameroo for output signals
  out_port_from_the_portconf_pio <= internal_out_port_from_the_portconf_pio;
  --vhdl renameroo for output signals
  out_port_from_the_status_led_pio <= internal_out_port_from_the_status_led_pio;
  --vhdl renameroo for output signals
  phasedone_from_the_altpll_0 <= internal_phasedone_from_the_altpll_0;
  --vhdl renameroo for output signals
  rTx_Dat_0_from_the_OpenMAC_0 <= internal_rTx_Dat_0_from_the_OpenMAC_0;
  --vhdl renameroo for output signals
  rTx_Dat_1_from_the_OpenMAC_0 <= internal_rTx_Dat_1_from_the_OpenMAC_0;
  --vhdl renameroo for output signals
  rTx_En_0_from_the_OpenMAC_0 <= internal_rTx_En_0_from_the_OpenMAC_0;
  --vhdl renameroo for output signals
  rTx_En_1_from_the_OpenMAC_0 <= internal_rTx_En_1_from_the_OpenMAC_0;
  --vhdl renameroo for output signals
  sce_from_the_epcs_flash_controller_0 <= internal_sce_from_the_epcs_flash_controller_0;
  --vhdl renameroo for output signals
  sdo_from_the_epcs_flash_controller_0 <= internal_sdo_from_the_epcs_flash_controller_0;
  --vhdl renameroo for output signals
  select_n_to_the_cfi_flash_0 <= internal_select_n_to_the_cfi_flash_0;
  --vhdl renameroo for output signals
  tri_state_bridge_0_address <= internal_tri_state_bridge_0_address;
  --vhdl renameroo for output signals
  tri_state_bridge_0_readn <= internal_tri_state_bridge_0_readn;
  --vhdl renameroo for output signals
  tri_state_bridge_0_writen <= internal_tri_state_bridge_0_writen;
  --vhdl renameroo for output signals
  zs_addr_from_the_sdram_0 <= internal_zs_addr_from_the_sdram_0;
  --vhdl renameroo for output signals
  zs_ba_from_the_sdram_0 <= internal_zs_ba_from_the_sdram_0;
  --vhdl renameroo for output signals
  zs_cas_n_from_the_sdram_0 <= internal_zs_cas_n_from_the_sdram_0;
  --vhdl renameroo for output signals
  zs_cke_from_the_sdram_0 <= internal_zs_cke_from_the_sdram_0;
  --vhdl renameroo for output signals
  zs_cs_n_from_the_sdram_0 <= internal_zs_cs_n_from_the_sdram_0;
  --vhdl renameroo for output signals
  zs_dqm_from_the_sdram_0 <= internal_zs_dqm_from_the_sdram_0;
  --vhdl renameroo for output signals
  zs_ras_n_from_the_sdram_0 <= internal_zs_ras_n_from_the_sdram_0;
  --vhdl renameroo for output signals
  zs_we_n_from_the_sdram_0 <= internal_zs_we_n_from_the_sdram_0;

end europa;


--synthesis translate_off

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity cfi_flash_0_lane0_module is 
        port (
              -- inputs:
                 signal data : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal rdaddress : IN STD_LOGIC_VECTOR (21 DOWNTO 0);
                 signal rdclken : IN STD_LOGIC;
                 signal wraddress : IN STD_LOGIC_VECTOR (21 DOWNTO 0);
                 signal wrclock : IN STD_LOGIC;
                 signal wren : IN STD_LOGIC;

              -- outputs:
                 signal q : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
              );
end entity cfi_flash_0_lane0_module;


architecture europa of cfi_flash_0_lane0_module is
              signal internal_q :  STD_LOGIC_VECTOR (7 DOWNTO 0);
              TYPE mem_array is ARRAY( 4194303 DOWNTO 0) of STD_LOGIC_VECTOR(7 DOWNTO 0);
              signal memory_has_been_read :  STD_LOGIC;
              signal read_address :  STD_LOGIC_VECTOR (21 DOWNTO 0);

      
FUNCTION convert_string_to_number(string_to_convert : STRING;
      final_char_index : NATURAL := 0)
RETURN NATURAL IS
   VARIABLE result: NATURAL := 0;
   VARIABLE current_index : NATURAL := 1;
   VARIABLE the_char : CHARACTER;

   BEGIN
      IF final_char_index = 0 THEN
         result := 0;
	 ELSE
         WHILE current_index <= final_char_index LOOP
            the_char := string_to_convert(current_index);
            IF    '0' <= the_char AND the_char <= '9' THEN
               result := result * 16 + character'pos(the_char) - character'pos('0');
            ELSIF 'A' <= the_char AND the_char <= 'F' THEN
               result := result * 16 + character'pos(the_char) - character'pos('A') + 10;
            ELSIF 'a' <= the_char AND the_char <= 'f' THEN
               result := result * 16 + character'pos(the_char) - character'pos('a') + 10;
            ELSE
               report "Ack, a formatting error!";
            END IF;
            current_index := current_index + 1;
         END LOOP;
      END IF; 
   RETURN result;
END convert_string_to_number;

 FUNCTION convert_string_to_std_logic(value : STRING; num_chars : INTEGER; mem_width_bits : INTEGER)
 RETURN STD_LOGIC_VECTOR is			   
     VARIABLE conv_string: std_logic_vector((mem_width_bits + 4)-1 downto 0);
     VARIABLE result : std_logic_vector((mem_width_bits -1) downto 0);
     VARIABLE curr_char : integer;
              
     BEGIN
     result := (others => '0');
     conv_string := (others => '0');
     
          FOR I IN 1 TO num_chars LOOP
	     curr_char := num_chars - (I-1);

             CASE value(I) IS
               WHEN '0' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0000";
               WHEN '1' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0001";
               WHEN '2' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0010";
               WHEN '3' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0011";
               WHEN '4' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0100";
               WHEN '5' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0101";
               WHEN '6' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0110";
               WHEN '7' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0111";
               WHEN '8' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1000";
               WHEN '9' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1001";
               WHEN 'A' | 'a' => conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1010";
               WHEN 'B' | 'b' => conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1011";
               WHEN 'C' | 'c' => conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1100";
               WHEN 'D' | 'd' => conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1101";
               WHEN 'E' | 'e' => conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1110";
               WHEN 'F' | 'f' => conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1111";
               WHEN 'X' | 'x' => conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "XXXX";
               WHEN ' ' => EXIT;
               WHEN HT  => exit;
               WHEN others =>
                  ASSERT False
                  REPORT "function From_Hex: string """ & value & """ contains non-hex character"
                       severity Error;
                  EXIT;
               END case;
            END loop;

          -- convert back to normal bit size
          result(mem_width_bits - 1 downto 0) := conv_string(mem_width_bits - 1 downto 0);

          RETURN result;
        END convert_string_to_std_logic;



begin
   process (wrclock, rdaddress) -- MG
    VARIABLE data_line : LINE;
    VARIABLE the_character_from_data_line : CHARACTER;
    VARIABLE b_munging_address : BOOLEAN := FALSE;
    VARIABLE converted_number : NATURAL := 0;
    VARIABLE found_string_array : STRING(1 TO 128);
    VARIABLE string_index : NATURAL := 0;
    VARIABLE line_length : NATURAL := 0;
    VARIABLE b_convert : BOOLEAN := FALSE;
    VARIABLE b_found_new_val : BOOLEAN := FALSE;
    VARIABLE load_address : NATURAL := 0;
    VARIABLE mem_index : NATURAL := 0;
    VARIABLE mem_init : BOOLEAN := FALSE;

    VARIABLE wr_address_internal : STD_LOGIC_VECTOR (21 DOWNTO 0) := (others => '0');
    FILE memory_contents_file : TEXT OPEN read_mode IS "cfi_flash_0_lane0.dat";  
    variable Marc_Gaucherons_Memory_Variable : mem_array; -- MG
    
    begin
   -- need an initialization process
   -- this process initializes the whole memory array from a named file by copying the
   -- contents of the *.dat file to the memory array.

   -- find the @<address> thingy to load the memory from this point 
IF(NOT mem_init) THEN
   WHILE NOT(endfile(memory_contents_file)) LOOP

      readline(memory_contents_file, data_line);
      line_length := data_line'LENGTH;


      WHILE line_length > 0 LOOP
         read(data_line, the_character_from_data_line);

	       -- check for the @ character indicating a new address wad
 	       -- if not found, we're either still reading the new address _or_loading data
         IF '@' = the_character_from_data_line AND NOT b_munging_address THEN
  	    b_munging_address := TRUE;
            b_found_new_val := TRUE; 
	    -- get the rest of characters before white space and then convert them
	    -- to a number
	 ELSE 

            IF (' ' = the_character_from_data_line AND b_found_new_val) 
		OR (line_length = 1) THEN
               b_convert := TRUE;
	    END IF;

            IF NOT(' ' = the_character_from_data_line) THEN
               string_index := string_index + 1;
               found_string_array(string_index) := the_character_from_data_line;
--               IF NOT(b_munging_address) THEN
--                 dat_string_array(string_index) := the_character_from_data_line;
--               END IF;
	       b_found_new_val := TRUE;
            END IF;
	 END IF;

     IF b_convert THEN

       IF b_munging_address THEN
          converted_number := convert_string_to_number(found_string_array, string_index);    
          load_address := converted_number;
          mem_index := load_address;
--          mem_index := load_address / 1;
          b_munging_address := FALSE;
       ELSE
	  IF (mem_index < 4194304) THEN
	    Marc_Gaucherons_Memory_Variable(mem_index) := convert_string_to_std_logic(found_string_array, string_index, 8);
            mem_index := mem_index + 1;
          END IF;
       END IF; 
       b_convert := FALSE;
       b_found_new_val := FALSE;
       string_index := 0;
    END IF;
    line_length := line_length - 1; 
    END LOOP;

END LOOP;
-- get the first _real_ block of data, sized to our memory width
-- and keep on loading.
  mem_init := TRUE;
END IF;
-- END OF READMEM



      -- Write data
      if wrclock'event and wrclock = '1' then
        wr_address_internal := wraddress;
        if wren = '1' then 
          Marc_Gaucherons_Memory_Variable(CONV_INTEGER(UNSIGNED(wr_address_internal))) := data;
        end if;
      end if;

      -- read data
      q <= Marc_Gaucherons_Memory_Variable(CONV_INTEGER(UNSIGNED(rdaddress)));
      


    end process;
end europa;

--synthesis translate_on


--synthesis read_comments_as_HDL on
--library altera;
--use altera.altera_europa_support_lib.all;
--
--library ieee;
--use ieee.std_logic_1164.all;
--use ieee.std_logic_arith.all;
--use ieee.std_logic_unsigned.all;
--
--library std;
--use std.textio.all;
--
--entity cfi_flash_0_lane0_module is 
--        port (
--              
--                 signal data : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
--                 signal rdaddress : IN STD_LOGIC_VECTOR (21 DOWNTO 0);
--                 signal rdclken : IN STD_LOGIC;
--                 signal wraddress : IN STD_LOGIC_VECTOR (21 DOWNTO 0);
--                 signal wrclock : IN STD_LOGIC;
--                 signal wren : IN STD_LOGIC;
--
--              
--                 signal q : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
--              );
--end entity cfi_flash_0_lane0_module;
--
--
--architecture europa of cfi_flash_0_lane0_module is
--  component lpm_ram_dp is
--GENERIC (
--      lpm_file : STRING;
--        lpm_hint : STRING;
--        lpm_indata : STRING;
--        lpm_outdata : STRING;
--        lpm_rdaddress_control : STRING;
--        lpm_width : NATURAL;
--        lpm_widthad : NATURAL;
--        lpm_wraddress_control : STRING;
--        suppress_memory_conversion_warnings : STRING
--      );
--    PORT (
--    signal q : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
--        signal rdaddress : IN STD_LOGIC_VECTOR (21 DOWNTO 0);
--        signal wren : IN STD_LOGIC;
--        signal wrclock : IN STD_LOGIC;
--        signal wraddress : IN STD_LOGIC_VECTOR (21 DOWNTO 0);
--        signal data : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
--        signal rdclken : IN STD_LOGIC
--      );
--  end component lpm_ram_dp;
--                signal internal_q :  STD_LOGIC_VECTOR (7 DOWNTO 0);
--                TYPE mem_array is ARRAY( 4194303 DOWNTO 0) of STD_LOGIC_VECTOR(7 DOWNTO 0);
--                signal memory_has_been_read :  STD_LOGIC;
--                signal read_address :  STD_LOGIC_VECTOR (21 DOWNTO 0);
--
--begin
--
--  process (rdaddress)
--  begin
--      read_address <= rdaddress;
--
--  end process;
--
--  lpm_ram_dp_component : lpm_ram_dp
--    generic map(
--      lpm_file => "cfi_flash_0_lane0.mif",
--      lpm_hint => "USE_EAB=ON",
--      lpm_indata => "REGISTERED",
--      lpm_outdata => "UNREGISTERED",
--      lpm_rdaddress_control => "UNREGISTERED",
--      lpm_width => 8,
--      lpm_widthad => 22,
--      lpm_wraddress_control => "REGISTERED",
--      suppress_memory_conversion_warnings => "ON"
--    )
--    port map(
--            data => data,
--            q => internal_q,
--            rdaddress => read_address,
--            rdclken => rdclken,
--            wraddress => wraddress,
--            wrclock => wrclock,
--            wren => wren
--    );
--
--  
--  q <= internal_q;
--end europa;
--
--synthesis read_comments_as_HDL off


-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 


--synthesis translate_off

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity cfi_flash_0_lane1_module is 
        port (
              -- inputs:
                 signal data : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal rdaddress : IN STD_LOGIC_VECTOR (21 DOWNTO 0);
                 signal rdclken : IN STD_LOGIC;
                 signal wraddress : IN STD_LOGIC_VECTOR (21 DOWNTO 0);
                 signal wrclock : IN STD_LOGIC;
                 signal wren : IN STD_LOGIC;

              -- outputs:
                 signal q : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
              );
end entity cfi_flash_0_lane1_module;


architecture europa of cfi_flash_0_lane1_module is
              signal internal_q1 :  STD_LOGIC_VECTOR (7 DOWNTO 0);
              TYPE mem_array is ARRAY( 4194303 DOWNTO 0) of STD_LOGIC_VECTOR(7 DOWNTO 0);
              signal memory_has_been_read :  STD_LOGIC;
              signal read_address :  STD_LOGIC_VECTOR (21 DOWNTO 0);

      
FUNCTION convert_string_to_number(string_to_convert : STRING;
      final_char_index : NATURAL := 0)
RETURN NATURAL IS
   VARIABLE result: NATURAL := 0;
   VARIABLE current_index : NATURAL := 1;
   VARIABLE the_char : CHARACTER;

   BEGIN
      IF final_char_index = 0 THEN
         result := 0;
	 ELSE
         WHILE current_index <= final_char_index LOOP
            the_char := string_to_convert(current_index);
            IF    '0' <= the_char AND the_char <= '9' THEN
               result := result * 16 + character'pos(the_char) - character'pos('0');
            ELSIF 'A' <= the_char AND the_char <= 'F' THEN
               result := result * 16 + character'pos(the_char) - character'pos('A') + 10;
            ELSIF 'a' <= the_char AND the_char <= 'f' THEN
               result := result * 16 + character'pos(the_char) - character'pos('a') + 10;
            ELSE
               report "Ack, a formatting error!";
            END IF;
            current_index := current_index + 1;
         END LOOP;
      END IF; 
   RETURN result;
END convert_string_to_number;

 FUNCTION convert_string_to_std_logic(value : STRING; num_chars : INTEGER; mem_width_bits : INTEGER)
 RETURN STD_LOGIC_VECTOR is			   
     VARIABLE conv_string: std_logic_vector((mem_width_bits + 4)-1 downto 0);
     VARIABLE result : std_logic_vector((mem_width_bits -1) downto 0);
     VARIABLE curr_char : integer;
              
     BEGIN
     result := (others => '0');
     conv_string := (others => '0');
     
          FOR I IN 1 TO num_chars LOOP
	     curr_char := num_chars - (I-1);

             CASE value(I) IS
               WHEN '0' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0000";
               WHEN '1' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0001";
               WHEN '2' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0010";
               WHEN '3' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0011";
               WHEN '4' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0100";
               WHEN '5' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0101";
               WHEN '6' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0110";
               WHEN '7' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0111";
               WHEN '8' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1000";
               WHEN '9' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1001";
               WHEN 'A' | 'a' => conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1010";
               WHEN 'B' | 'b' => conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1011";
               WHEN 'C' | 'c' => conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1100";
               WHEN 'D' | 'd' => conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1101";
               WHEN 'E' | 'e' => conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1110";
               WHEN 'F' | 'f' => conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1111";
               WHEN 'X' | 'x' => conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "XXXX";
               WHEN ' ' => EXIT;
               WHEN HT  => exit;
               WHEN others =>
                  ASSERT False
                  REPORT "function From_Hex: string """ & value & """ contains non-hex character"
                       severity Error;
                  EXIT;
               END case;
            END loop;

          -- convert back to normal bit size
          result(mem_width_bits - 1 downto 0) := conv_string(mem_width_bits - 1 downto 0);

          RETURN result;
        END convert_string_to_std_logic;



begin
   process (wrclock, rdaddress) -- MG
    VARIABLE data_line : LINE;
    VARIABLE the_character_from_data_line : CHARACTER;
    VARIABLE b_munging_address : BOOLEAN := FALSE;
    VARIABLE converted_number : NATURAL := 0;
    VARIABLE found_string_array : STRING(1 TO 128);
    VARIABLE string_index : NATURAL := 0;
    VARIABLE line_length : NATURAL := 0;
    VARIABLE b_convert : BOOLEAN := FALSE;
    VARIABLE b_found_new_val : BOOLEAN := FALSE;
    VARIABLE load_address : NATURAL := 0;
    VARIABLE mem_index : NATURAL := 0;
    VARIABLE mem_init : BOOLEAN := FALSE;

    VARIABLE wr_address_internal : STD_LOGIC_VECTOR (21 DOWNTO 0) := (others => '0');
    FILE memory_contents_file : TEXT OPEN read_mode IS "cfi_flash_0_lane1.dat";  
    variable Marc_Gaucherons_Memory_Variable : mem_array; -- MG
    
    begin
   -- need an initialization process
   -- this process initializes the whole memory array from a named file by copying the
   -- contents of the *.dat file to the memory array.

   -- find the @<address> thingy to load the memory from this point 
IF(NOT mem_init) THEN
   WHILE NOT(endfile(memory_contents_file)) LOOP

      readline(memory_contents_file, data_line);
      line_length := data_line'LENGTH;


      WHILE line_length > 0 LOOP
         read(data_line, the_character_from_data_line);

	       -- check for the @ character indicating a new address wad
 	       -- if not found, we're either still reading the new address _or_loading data
         IF '@' = the_character_from_data_line AND NOT b_munging_address THEN
  	    b_munging_address := TRUE;
            b_found_new_val := TRUE; 
	    -- get the rest of characters before white space and then convert them
	    -- to a number
	 ELSE 

            IF (' ' = the_character_from_data_line AND b_found_new_val) 
		OR (line_length = 1) THEN
               b_convert := TRUE;
	    END IF;

            IF NOT(' ' = the_character_from_data_line) THEN
               string_index := string_index + 1;
               found_string_array(string_index) := the_character_from_data_line;
--               IF NOT(b_munging_address) THEN
--                 dat_string_array(string_index) := the_character_from_data_line;
--               END IF;
	       b_found_new_val := TRUE;
            END IF;
	 END IF;

     IF b_convert THEN

       IF b_munging_address THEN
          converted_number := convert_string_to_number(found_string_array, string_index);    
          load_address := converted_number;
          mem_index := load_address;
--          mem_index := load_address / 1;
          b_munging_address := FALSE;
       ELSE
	  IF (mem_index < 4194304) THEN
	    Marc_Gaucherons_Memory_Variable(mem_index) := convert_string_to_std_logic(found_string_array, string_index, 8);
            mem_index := mem_index + 1;
          END IF;
       END IF; 
       b_convert := FALSE;
       b_found_new_val := FALSE;
       string_index := 0;
    END IF;
    line_length := line_length - 1; 
    END LOOP;

END LOOP;
-- get the first _real_ block of data, sized to our memory width
-- and keep on loading.
  mem_init := TRUE;
END IF;
-- END OF READMEM



      -- Write data
      if wrclock'event and wrclock = '1' then
        wr_address_internal := wraddress;
        if wren = '1' then 
          Marc_Gaucherons_Memory_Variable(CONV_INTEGER(UNSIGNED(wr_address_internal))) := data;
        end if;
      end if;

      -- read data
      q <= Marc_Gaucherons_Memory_Variable(CONV_INTEGER(UNSIGNED(rdaddress)));
      


    end process;
end europa;

--synthesis translate_on


--synthesis read_comments_as_HDL on
--library altera;
--use altera.altera_europa_support_lib.all;
--
--library ieee;
--use ieee.std_logic_1164.all;
--use ieee.std_logic_arith.all;
--use ieee.std_logic_unsigned.all;
--
--library std;
--use std.textio.all;
--
--entity cfi_flash_0_lane1_module is 
--        port (
--              
--                 signal data : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
--                 signal rdaddress : IN STD_LOGIC_VECTOR (21 DOWNTO 0);
--                 signal rdclken : IN STD_LOGIC;
--                 signal wraddress : IN STD_LOGIC_VECTOR (21 DOWNTO 0);
--                 signal wrclock : IN STD_LOGIC;
--                 signal wren : IN STD_LOGIC;
--
--              
--                 signal q : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
--              );
--end entity cfi_flash_0_lane1_module;
--
--
--architecture europa of cfi_flash_0_lane1_module is
--  component lpm_ram_dp is
--GENERIC (
--      lpm_file : STRING;
--        lpm_hint : STRING;
--        lpm_indata : STRING;
--        lpm_outdata : STRING;
--        lpm_rdaddress_control : STRING;
--        lpm_width : NATURAL;
--        lpm_widthad : NATURAL;
--        lpm_wraddress_control : STRING;
--        suppress_memory_conversion_warnings : STRING
--      );
--    PORT (
--    signal q : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
--        signal rdaddress : IN STD_LOGIC_VECTOR (21 DOWNTO 0);
--        signal wren : IN STD_LOGIC;
--        signal wrclock : IN STD_LOGIC;
--        signal wraddress : IN STD_LOGIC_VECTOR (21 DOWNTO 0);
--        signal data : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
--        signal rdclken : IN STD_LOGIC
--      );
--  end component lpm_ram_dp;
--                signal internal_q1 :  STD_LOGIC_VECTOR (7 DOWNTO 0);
--                TYPE mem_array is ARRAY( 4194303 DOWNTO 0) of STD_LOGIC_VECTOR(7 DOWNTO 0);
--                signal memory_has_been_read :  STD_LOGIC;
--                signal read_address :  STD_LOGIC_VECTOR (21 DOWNTO 0);
--
--begin
--
--  process (rdaddress)
--  begin
--      read_address <= rdaddress;
--
--  end process;
--
--  lpm_ram_dp_component : lpm_ram_dp
--    generic map(
--      lpm_file => "cfi_flash_0_lane1.mif",
--      lpm_hint => "USE_EAB=ON",
--      lpm_indata => "REGISTERED",
--      lpm_outdata => "UNREGISTERED",
--      lpm_rdaddress_control => "UNREGISTERED",
--      lpm_width => 8,
--      lpm_widthad => 22,
--      lpm_wraddress_control => "REGISTERED",
--      suppress_memory_conversion_warnings => "ON"
--    )
--    port map(
--            data => data,
--            q => internal_q1,
--            rdaddress => read_address,
--            rdclken => rdclken,
--            wraddress => wraddress,
--            wrclock => wrclock,
--            wren => wren
--    );
--
--  
--  q <= internal_q1;
--end europa;
--
--synthesis read_comments_as_HDL off


-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity cfi_flash_0 is 
        port (
              -- inputs:
                 signal address : IN STD_LOGIC_VECTOR (21 DOWNTO 0);
                 signal read_n : IN STD_LOGIC;
                 signal select_n : IN STD_LOGIC;
                 signal write_n : IN STD_LOGIC;

              -- outputs:
                 signal data : INOUT STD_LOGIC_VECTOR (15 DOWNTO 0)
              );
end entity cfi_flash_0;


architecture europa of cfi_flash_0 is
--synthesis translate_off
component cfi_flash_0_lane0_module is 
           port (
                 -- inputs:
                    signal data : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal rdaddress : IN STD_LOGIC_VECTOR (21 DOWNTO 0);
                    signal rdclken : IN STD_LOGIC;
                    signal wraddress : IN STD_LOGIC_VECTOR (21 DOWNTO 0);
                    signal wrclock : IN STD_LOGIC;
                    signal wren : IN STD_LOGIC;

                 -- outputs:
                    signal q : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
                 );
end component cfi_flash_0_lane0_module;

component cfi_flash_0_lane1_module is 
           port (
                 -- inputs:
                    signal data : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal rdaddress : IN STD_LOGIC_VECTOR (21 DOWNTO 0);
                    signal rdclken : IN STD_LOGIC;
                    signal wraddress : IN STD_LOGIC_VECTOR (21 DOWNTO 0);
                    signal wrclock : IN STD_LOGIC;
                    signal wren : IN STD_LOGIC;

                 -- outputs:
                    signal q : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
                 );
end component cfi_flash_0_lane1_module;

--synthesis translate_on
                signal data_0 :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal data_1 :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal logic_vector_gasket :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal module_input16 :  STD_LOGIC;
                signal module_input17 :  STD_LOGIC;
                signal module_input18 :  STD_LOGIC;
                signal module_input19 :  STD_LOGIC;
                signal q_0 :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal q_1 :  STD_LOGIC_VECTOR (7 DOWNTO 0);

begin

  --s1, which is an e_ptf_slave
--synthesis translate_off
    logic_vector_gasket <= data;
    data_0 <= logic_vector_gasket(7 DOWNTO 0);
    --cfi_flash_0_lane0, which is an e_ram
    cfi_flash_0_lane0 : cfi_flash_0_lane0_module
      port map(
        q => q_0,
        data => data_0,
        rdaddress => address,
        rdclken => module_input16,
        wraddress => address,
        wrclock => write_n,
        wren => module_input17
      );

    module_input16 <= std_logic'('1');
    module_input17 <= NOT select_n;

    data_1 <= logic_vector_gasket(15 DOWNTO 8);
    --cfi_flash_0_lane1, which is an e_ram
    cfi_flash_0_lane1 : cfi_flash_0_lane1_module
      port map(
        q => q_1,
        data => data_1,
        rdaddress => address,
        rdclken => module_input18,
        wraddress => address,
        wrclock => write_n,
        wren => module_input19
      );

    module_input18 <= std_logic'('1');
    module_input19 <= NOT select_n;

    data <= A_WE_StdLogicVector((std_logic'(((NOT select_n AND NOT read_n))) = '1'), (q_1 & q_0), A_REP(std_logic'('Z'), 16));
--synthesis translate_on

end europa;


--synthesis translate_off

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;



-- <ALTERA_NOTE> CODE INSERTED BETWEEN HERE
--add your libraries here
-- AND HERE WILL BE PRESERVED </ALTERA_NOTE>

entity test_bench is 
end entity test_bench;


architecture europa of test_bench is
component niosII_openMac is 
           port (
                 -- 1) global signals:
                    signal clk100Meg180 : OUT STD_LOGIC;
                    signal clk25Meg : OUT STD_LOGIC;
                    signal clk50Meg : OUT STD_LOGIC;
                    signal clk90Meg : OUT STD_LOGIC;
                    signal clk90MegSDRAM : OUT STD_LOGIC;
                    signal clk_0 : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- the_OpenMAC_0
                    signal mii_Clk_from_the_OpenMAC_0 : OUT STD_LOGIC;
                    signal mii_Di_to_the_OpenMAC_0 : IN STD_LOGIC;
                    signal mii_Do_from_the_OpenMAC_0 : OUT STD_LOGIC;
                    signal mii_Doe_from_the_OpenMAC_0 : OUT STD_LOGIC;
                    signal mii_nResetOut_from_the_OpenMAC_0 : OUT STD_LOGIC;
                    signal rCrs_Dv_0_to_the_OpenMAC_0 : IN STD_LOGIC;
                    signal rCrs_Dv_1_to_the_OpenMAC_0 : IN STD_LOGIC;
                    signal rRx_Dat_0_to_the_OpenMAC_0 : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal rRx_Dat_1_to_the_OpenMAC_0 : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal rTx_Dat_0_from_the_OpenMAC_0 : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal rTx_Dat_1_from_the_OpenMAC_0 : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal rTx_En_0_from_the_OpenMAC_0 : OUT STD_LOGIC;
                    signal rTx_En_1_from_the_OpenMAC_0 : OUT STD_LOGIC;

                 -- the_altpll_0
                    signal locked_from_the_altpll_0 : OUT STD_LOGIC;
                    signal phasedone_from_the_altpll_0 : OUT STD_LOGIC;

                 -- the_button_pio
                    signal in_port_to_the_button_pio : IN STD_LOGIC_VECTOR (7 DOWNTO 0);

                 -- the_digio_pio
                    signal bidir_port_to_and_from_the_digio_pio : INOUT STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- the_epcs_flash_controller_0
                    signal data0_to_the_epcs_flash_controller_0 : IN STD_LOGIC;
                    signal dclk_from_the_epcs_flash_controller_0 : OUT STD_LOGIC;
                    signal sce_from_the_epcs_flash_controller_0 : OUT STD_LOGIC;
                    signal sdo_from_the_epcs_flash_controller_0 : OUT STD_LOGIC;

                 -- the_irq_gen
                    signal out_port_from_the_irq_gen : OUT STD_LOGIC;

                 -- the_node_switch_pio
                    signal in_port_to_the_node_switch_pio : IN STD_LOGIC_VECTOR (7 DOWNTO 0);

                 -- the_portconf_pio
                    signal in_port_to_the_portconf_pio : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal out_port_from_the_portconf_pio : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);

                 -- the_sdram_0
                    signal zs_addr_from_the_sdram_0 : OUT STD_LOGIC_VECTOR (11 DOWNTO 0);
                    signal zs_ba_from_the_sdram_0 : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal zs_cas_n_from_the_sdram_0 : OUT STD_LOGIC;
                    signal zs_cke_from_the_sdram_0 : OUT STD_LOGIC;
                    signal zs_cs_n_from_the_sdram_0 : OUT STD_LOGIC;
                    signal zs_dq_to_and_from_the_sdram_0 : INOUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal zs_dqm_from_the_sdram_0 : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal zs_ras_n_from_the_sdram_0 : OUT STD_LOGIC;
                    signal zs_we_n_from_the_sdram_0 : OUT STD_LOGIC;

                 -- the_status_led_pio
                    signal out_port_from_the_status_led_pio : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);

                 -- the_sync_irq
                    signal in_port_to_the_sync_irq : IN STD_LOGIC;

                 -- the_tri_state_bridge_0_avalon_slave
                    signal ben_to_the_DBC3C40_SRAM_0 : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal ncs_to_the_DBC3C40_SRAM_0 : OUT STD_LOGIC;
                    signal select_n_to_the_cfi_flash_0 : OUT STD_LOGIC;
                    signal tri_state_bridge_0_address : OUT STD_LOGIC_VECTOR (22 DOWNTO 0);
                    signal tri_state_bridge_0_data : INOUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal tri_state_bridge_0_readn : OUT STD_LOGIC;
                    signal tri_state_bridge_0_writen : OUT STD_LOGIC
                 );
end component niosII_openMac;

component cfi_flash_0 is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (21 DOWNTO 0);
                    signal read_n : IN STD_LOGIC;
                    signal select_n : IN STD_LOGIC;
                    signal write_n : IN STD_LOGIC;

                 -- outputs:
                    signal data : INOUT STD_LOGIC_VECTOR (15 DOWNTO 0)
                 );
end component cfi_flash_0;

component sdram_0_test_component is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal zs_addr : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
                    signal zs_ba : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal zs_cas_n : IN STD_LOGIC;
                    signal zs_cke : IN STD_LOGIC;
                    signal zs_cs_n : IN STD_LOGIC;
                    signal zs_dqm : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal zs_ras_n : IN STD_LOGIC;
                    signal zs_we_n : IN STD_LOGIC;

                 -- outputs:
                    signal zs_dq : INOUT STD_LOGIC_VECTOR (31 DOWNTO 0)
                 );
end component sdram_0_test_component;

                signal ben_to_the_DBC3C40_SRAM_0 :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal bidir_port_to_and_from_the_digio_pio :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal clk :  STD_LOGIC;
                signal clk100Meg180 :  STD_LOGIC;
                signal clk25Meg :  STD_LOGIC;
                signal clk50Meg :  STD_LOGIC;
                signal clk90Meg :  STD_LOGIC;
                signal clk90MegSDRAM :  STD_LOGIC;
                signal clk_0 :  STD_LOGIC;
                signal clock_crossing_0_m1_endofpacket :  STD_LOGIC;
                signal clock_crossing_0_s1_endofpacket_from_sa :  STD_LOGIC;
                signal clock_crossing_1_m1_endofpacket :  STD_LOGIC;
                signal clock_crossing_1_s1_endofpacket_from_sa :  STD_LOGIC;
                signal data0_to_the_epcs_flash_controller_0 :  STD_LOGIC;
                signal dclk_from_the_epcs_flash_controller_0 :  STD_LOGIC;
                signal epcs_flash_controller_0_epcs_control_port_dataavailable_from_sa :  STD_LOGIC;
                signal epcs_flash_controller_0_epcs_control_port_endofpacket_from_sa :  STD_LOGIC;
                signal epcs_flash_controller_0_epcs_control_port_readyfordata_from_sa :  STD_LOGIC;
                signal in_port_to_the_button_pio :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal in_port_to_the_node_switch_pio :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal in_port_to_the_portconf_pio :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal in_port_to_the_sync_irq :  STD_LOGIC;
                signal jtag_uart_0_avalon_jtag_slave_dataavailable_from_sa :  STD_LOGIC;
                signal jtag_uart_0_avalon_jtag_slave_readyfordata_from_sa :  STD_LOGIC;
                signal jtag_uart_1_avalon_jtag_slave_dataavailable_from_sa :  STD_LOGIC;
                signal jtag_uart_1_avalon_jtag_slave_readyfordata_from_sa :  STD_LOGIC;
                signal locked_from_the_altpll_0 :  STD_LOGIC;
                signal mii_Clk_from_the_OpenMAC_0 :  STD_LOGIC;
                signal mii_Di_to_the_OpenMAC_0 :  STD_LOGIC;
                signal mii_Do_from_the_OpenMAC_0 :  STD_LOGIC;
                signal mii_Doe_from_the_OpenMAC_0 :  STD_LOGIC;
                signal mii_nResetOut_from_the_OpenMAC_0 :  STD_LOGIC;
                signal module_input20 :  STD_LOGIC_VECTOR (21 DOWNTO 0);
                signal ncs_to_the_DBC3C40_SRAM_0 :  STD_LOGIC;
                signal niosII_openMac_clock_0_in_endofpacket_from_sa :  STD_LOGIC;
                signal niosII_openMac_clock_0_out_endofpacket :  STD_LOGIC;
                signal niosII_openMac_clock_1_in_endofpacket_from_sa :  STD_LOGIC;
                signal niosII_openMac_clock_1_out_endofpacket :  STD_LOGIC;
                signal niosII_openMac_clock_1_out_nativeaddress :  STD_LOGIC;
                signal niosII_openMac_clock_2_in_endofpacket_from_sa :  STD_LOGIC;
                signal niosII_openMac_clock_2_out_endofpacket :  STD_LOGIC;
                signal niosII_openMac_clock_2_out_nativeaddress :  STD_LOGIC_VECTOR (11 DOWNTO 0);
                signal niosII_openMac_clock_3_in_endofpacket_from_sa :  STD_LOGIC;
                signal niosII_openMac_clock_3_out_endofpacket :  STD_LOGIC;
                signal niosII_openMac_clock_3_out_nativeaddress :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal niosII_openMac_clock_4_in_endofpacket_from_sa :  STD_LOGIC;
                signal niosII_openMac_clock_4_out_endofpacket :  STD_LOGIC;
                signal out_port_from_the_irq_gen :  STD_LOGIC;
                signal out_port_from_the_portconf_pio :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal out_port_from_the_status_led_pio :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal phasedone_from_the_altpll_0 :  STD_LOGIC;
                signal rCrs_Dv_0_to_the_OpenMAC_0 :  STD_LOGIC;
                signal rCrs_Dv_1_to_the_OpenMAC_0 :  STD_LOGIC;
                signal rRx_Dat_0_to_the_OpenMAC_0 :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal rRx_Dat_1_to_the_OpenMAC_0 :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal rTx_Dat_0_from_the_OpenMAC_0 :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal rTx_Dat_1_from_the_OpenMAC_0 :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal rTx_En_0_from_the_OpenMAC_0 :  STD_LOGIC;
                signal rTx_En_1_from_the_OpenMAC_0 :  STD_LOGIC;
                signal reset_n :  STD_LOGIC;
                signal sce_from_the_epcs_flash_controller_0 :  STD_LOGIC;
                signal sdo_from_the_epcs_flash_controller_0 :  STD_LOGIC;
                signal select_n_to_the_cfi_flash_0 :  STD_LOGIC;
                signal tri_state_bridge_0_address :  STD_LOGIC_VECTOR (22 DOWNTO 0);
                signal tri_state_bridge_0_data :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal tri_state_bridge_0_readn :  STD_LOGIC;
                signal tri_state_bridge_0_writen :  STD_LOGIC;
                signal zs_addr_from_the_sdram_0 :  STD_LOGIC_VECTOR (11 DOWNTO 0);
                signal zs_ba_from_the_sdram_0 :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal zs_cas_n_from_the_sdram_0 :  STD_LOGIC;
                signal zs_cke_from_the_sdram_0 :  STD_LOGIC;
                signal zs_cs_n_from_the_sdram_0 :  STD_LOGIC;
                signal zs_dq_to_and_from_the_sdram_0 :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal zs_dqm_from_the_sdram_0 :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal zs_ras_n_from_the_sdram_0 :  STD_LOGIC;
                signal zs_we_n_from_the_sdram_0 :  STD_LOGIC;


-- <ALTERA_NOTE> CODE INSERTED BETWEEN HERE
--add your component and signal declaration here
-- AND HERE WILL BE PRESERVED </ALTERA_NOTE>


begin

  --Set us up the Dut
  DUT : niosII_openMac
    port map(
      ben_to_the_DBC3C40_SRAM_0 => ben_to_the_DBC3C40_SRAM_0,
      bidir_port_to_and_from_the_digio_pio => bidir_port_to_and_from_the_digio_pio,
      clk100Meg180 => clk100Meg180,
      clk25Meg => clk25Meg,
      clk50Meg => clk50Meg,
      clk90Meg => clk90Meg,
      clk90MegSDRAM => clk90MegSDRAM,
      dclk_from_the_epcs_flash_controller_0 => dclk_from_the_epcs_flash_controller_0,
      locked_from_the_altpll_0 => locked_from_the_altpll_0,
      mii_Clk_from_the_OpenMAC_0 => mii_Clk_from_the_OpenMAC_0,
      mii_Do_from_the_OpenMAC_0 => mii_Do_from_the_OpenMAC_0,
      mii_Doe_from_the_OpenMAC_0 => mii_Doe_from_the_OpenMAC_0,
      mii_nResetOut_from_the_OpenMAC_0 => mii_nResetOut_from_the_OpenMAC_0,
      ncs_to_the_DBC3C40_SRAM_0 => ncs_to_the_DBC3C40_SRAM_0,
      out_port_from_the_irq_gen => out_port_from_the_irq_gen,
      out_port_from_the_portconf_pio => out_port_from_the_portconf_pio,
      out_port_from_the_status_led_pio => out_port_from_the_status_led_pio,
      phasedone_from_the_altpll_0 => phasedone_from_the_altpll_0,
      rTx_Dat_0_from_the_OpenMAC_0 => rTx_Dat_0_from_the_OpenMAC_0,
      rTx_Dat_1_from_the_OpenMAC_0 => rTx_Dat_1_from_the_OpenMAC_0,
      rTx_En_0_from_the_OpenMAC_0 => rTx_En_0_from_the_OpenMAC_0,
      rTx_En_1_from_the_OpenMAC_0 => rTx_En_1_from_the_OpenMAC_0,
      sce_from_the_epcs_flash_controller_0 => sce_from_the_epcs_flash_controller_0,
      sdo_from_the_epcs_flash_controller_0 => sdo_from_the_epcs_flash_controller_0,
      select_n_to_the_cfi_flash_0 => select_n_to_the_cfi_flash_0,
      tri_state_bridge_0_address => tri_state_bridge_0_address,
      tri_state_bridge_0_data => tri_state_bridge_0_data,
      tri_state_bridge_0_readn => tri_state_bridge_0_readn,
      tri_state_bridge_0_writen => tri_state_bridge_0_writen,
      zs_addr_from_the_sdram_0 => zs_addr_from_the_sdram_0,
      zs_ba_from_the_sdram_0 => zs_ba_from_the_sdram_0,
      zs_cas_n_from_the_sdram_0 => zs_cas_n_from_the_sdram_0,
      zs_cke_from_the_sdram_0 => zs_cke_from_the_sdram_0,
      zs_cs_n_from_the_sdram_0 => zs_cs_n_from_the_sdram_0,
      zs_dq_to_and_from_the_sdram_0 => zs_dq_to_and_from_the_sdram_0,
      zs_dqm_from_the_sdram_0 => zs_dqm_from_the_sdram_0,
      zs_ras_n_from_the_sdram_0 => zs_ras_n_from_the_sdram_0,
      zs_we_n_from_the_sdram_0 => zs_we_n_from_the_sdram_0,
      clk_0 => clk_0,
      data0_to_the_epcs_flash_controller_0 => data0_to_the_epcs_flash_controller_0,
      in_port_to_the_button_pio => in_port_to_the_button_pio,
      in_port_to_the_node_switch_pio => in_port_to_the_node_switch_pio,
      in_port_to_the_portconf_pio => in_port_to_the_portconf_pio,
      in_port_to_the_sync_irq => in_port_to_the_sync_irq,
      mii_Di_to_the_OpenMAC_0 => mii_Di_to_the_OpenMAC_0,
      rCrs_Dv_0_to_the_OpenMAC_0 => rCrs_Dv_0_to_the_OpenMAC_0,
      rCrs_Dv_1_to_the_OpenMAC_0 => rCrs_Dv_1_to_the_OpenMAC_0,
      rRx_Dat_0_to_the_OpenMAC_0 => rRx_Dat_0_to_the_OpenMAC_0,
      rRx_Dat_1_to_the_OpenMAC_0 => rRx_Dat_1_to_the_OpenMAC_0,
      reset_n => reset_n
    );


  --the_cfi_flash_0, which is an e_ptf_instance
  the_cfi_flash_0 : cfi_flash_0
    port map(
      data => tri_state_bridge_0_data,
      address => module_input20,
      read_n => tri_state_bridge_0_readn,
      select_n => select_n_to_the_cfi_flash_0,
      write_n => tri_state_bridge_0_writen
    );

  module_input20 <= tri_state_bridge_0_address(22 DOWNTO 1);

  --the_sdram_0_test_component, which is an e_instance
  the_sdram_0_test_component : sdram_0_test_component
    port map(
      zs_dq => zs_dq_to_and_from_the_sdram_0,
      clk => clk90Meg,
      zs_addr => zs_addr_from_the_sdram_0,
      zs_ba => zs_ba_from_the_sdram_0,
      zs_cas_n => zs_cas_n_from_the_sdram_0,
      zs_cke => zs_cke_from_the_sdram_0,
      zs_cs_n => zs_cs_n_from_the_sdram_0,
      zs_dqm => zs_dqm_from_the_sdram_0,
      zs_ras_n => zs_ras_n_from_the_sdram_0,
      zs_we_n => zs_we_n_from_the_sdram_0
    );


  process
  begin
    clk_0 <= '0';
    loop
       wait for 10 ns;
       clk_0 <= not clk_0;
    end loop;
  end process;
  PROCESS
    BEGIN
       reset_n <= '0';
       wait for 200 ns;
       reset_n <= '1'; 
    WAIT;
  END PROCESS;


-- <ALTERA_NOTE> CODE INSERTED BETWEEN HERE
--add additional architecture here
-- AND HERE WILL BE PRESERVED </ALTERA_NOTE>


end europa;



--synthesis translate_on
